-- srec2vhdl table generator
-- for input file hex_display.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"93874186",
           5 => x"13874186",
           6 => x"63e4e702",
           7 => x"b7070020",
           8 => x"1307401f",
           9 => x"93870700",
          10 => x"93864186",
          11 => x"63e2d702",
          12 => x"ef00c00e",
          13 => x"ef004005",
          14 => x"13050000",
          15 => x"ef00400a",
          16 => x"23a00700",
          17 => x"83a60700",
          18 => x"93874700",
          19 => x"6ff0dffc",
          20 => x"03260700",
          21 => x"93874700",
          22 => x"13074700",
          23 => x"23aec7fe",
          24 => x"6ff0dffc",
          25 => x"13030500",
          26 => x"630e0600",
          27 => x"83830500",
          28 => x"23007300",
          29 => x"1306f6ff",
          30 => x"13031300",
          31 => x"93851500",
          32 => x"e31606fe",
          33 => x"67800000",
          34 => x"130101fe",
          35 => x"13060001",
          36 => x"9305001e",
          37 => x"13050100",
          38 => x"232e1100",
          39 => x"eff09ffc",
          40 => x"b70600f0",
          41 => x"83a70600",
          42 => x"13d74700",
          43 => x"1377f700",
          44 => x"93f7f700",
          45 => x"13070701",
          46 => x"93870701",
          47 => x"33072700",
          48 => x"b3872700",
          49 => x"034707ff",
          50 => x"83c707ff",
          51 => x"13178701",
          52 => x"93970701",
          53 => x"b367f700",
          54 => x"23a2f600",
          55 => x"6ff09ffc",
          56 => x"130101ff",
          57 => x"23248100",
          58 => x"23261100",
          59 => x"93070000",
          60 => x"13040500",
          61 => x"63880700",
          62 => x"93050000",
          63 => x"97000000",
          64 => x"e7000000",
          65 => x"0325001f",
          66 => x"83278502",
          67 => x"63840700",
          68 => x"e7800700",
          69 => x"13050400",
          70 => x"ef000009",
          71 => x"130101ff",
          72 => x"23248100",
          73 => x"23229100",
          74 => x"9307401f",
          75 => x"1304401f",
          76 => x"3304f440",
          77 => x"23202101",
          78 => x"23261100",
          79 => x"13542440",
          80 => x"9304401f",
          81 => x"13090000",
          82 => x"631c8902",
          83 => x"9307401f",
          84 => x"1304401f",
          85 => x"3304f440",
          86 => x"13542440",
          87 => x"9304401f",
          88 => x"13090000",
          89 => x"63188902",
          90 => x"8320c100",
          91 => x"03248100",
          92 => x"83244100",
          93 => x"03290100",
          94 => x"13010101",
          95 => x"67800000",
          96 => x"83a70400",
          97 => x"13091900",
          98 => x"93844400",
          99 => x"e7800700",
         100 => x"6ff09ffb",
         101 => x"83a70400",
         102 => x"13091900",
         103 => x"93844400",
         104 => x"e7800700",
         105 => x"6ff01ffc",
         106 => x"9308d005",
         107 => x"73000000",
         108 => x"63520502",
         109 => x"130101ff",
         110 => x"23248100",
         111 => x"13040500",
         112 => x"23261100",
         113 => x"33048040",
         114 => x"ef000001",
         115 => x"23208500",
         116 => x"6f000000",
         117 => x"6f000000",
         118 => x"03a50186",
         119 => x"67800000",
         120 => x"40792430",
         121 => x"19120278",
         122 => x"00100803",
         123 => x"4621060e",
         124 => x"00000020",
         125 => x"00000000",
         126 => x"00000000",
         127 => x"00000000",
         128 => x"00000000",
         129 => x"00000000",
         130 => x"00000000",
         131 => x"00000000",
         132 => x"00000000",
         133 => x"00000000",
         134 => x"00000000",
         135 => x"00000000",
         136 => x"00000000",
         137 => x"00000000",
         138 => x"00000000",
         139 => x"00000000",
         140 => x"00000000",
         141 => x"00000000",
         142 => x"00000000",
         143 => x"00000000",
         144 => x"00000000",
         145 => x"00000000",
         146 => x"00000000",
         147 => x"00000000",
         148 => x"00000000",
         149 => x"00000020",
        others => (others => '-')
    );
end package processor_common_rom;
