-- srec2vhdl table generator
-- for input file shift.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97",    1 => x"11",    2 => x"00",    3 => x"20", 
           4 => x"93",    5 => x"81",    6 => x"01",    7 => x"80", 
           8 => x"17",    9 => x"41",   10 => x"00",   11 => x"20", 
          12 => x"13",   13 => x"01",   14 => x"81",   15 => x"ff", 
          16 => x"97",   17 => x"00",   18 => x"00",   19 => x"00", 
          20 => x"e7",   21 => x"80",   22 => x"c0",   23 => x"00", 
          24 => x"6f",   25 => x"00",   26 => x"00",   27 => x"00", 
          28 => x"13",   29 => x"01",   30 => x"01",   31 => x"fe", 
          32 => x"23",   33 => x"2e",   34 => x"81",   35 => x"00", 
          36 => x"13",   37 => x"04",   38 => x"01",   39 => x"02", 
          40 => x"93",   41 => x"07",   42 => x"10",   43 => x"00", 
          44 => x"23",   45 => x"26",   46 => x"f4",   47 => x"fe", 
          48 => x"83",   49 => x"27",   50 => x"c4",   51 => x"fe", 
          52 => x"93",   53 => x"97",   54 => x"47",   55 => x"00", 
          56 => x"23",   57 => x"26",   58 => x"f4",   59 => x"fe", 
          60 => x"93",   61 => x"07",   62 => x"00",   63 => x"00", 
          64 => x"13",   65 => x"85",   66 => x"07",   67 => x"00", 
          68 => x"03",   69 => x"24",   70 => x"c1",   71 => x"01", 
          72 => x"13",   73 => x"01",   74 => x"01",   75 => x"02", 
          76 => x"67",   77 => x"80",   78 => x"00",   79 => x"00", 
        others => (others => '-')
    );
end package processor_common_rom;
