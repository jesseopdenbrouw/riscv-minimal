-- srec2vhdl table generator
-- for input file exp.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"1387c186",
           5 => x"9386c186",
           6 => x"637ed700",
           7 => x"9387c186",
           8 => x"23800700",
           9 => x"13870700",
          10 => x"03470700",
          11 => x"93871700",
          12 => x"e398d7fe",
          13 => x"b7070020",
          14 => x"13870700",
          15 => x"1386c186",
          16 => x"6374c702",
          17 => x"b7160000",
          18 => x"9386060b",
          19 => x"93870700",
          20 => x"03c70600",
          21 => x"93871700",
          22 => x"93861600",
          23 => x"1377f70f",
          24 => x"a38fe7fe",
          25 => x"e396c7fe",
          26 => x"ef001063",
          27 => x"ef009059",
          28 => x"ef00506c",
          29 => x"37078000",
          30 => x"130101ff",
          31 => x"1307f7ff",
          32 => x"b377a700",
          33 => x"23248100",
          34 => x"23229100",
          35 => x"13547501",
          36 => x"9354f501",
          37 => x"13d57501",
          38 => x"3377b700",
          39 => x"1374f40f",
          40 => x"1375f50f",
          41 => x"23261100",
          42 => x"23202101",
          43 => x"93d5f501",
          44 => x"93973700",
          45 => x"13173700",
          46 => x"b306a440",
          47 => x"6396b418",
          48 => x"6358d00a",
          49 => x"63100504",
          50 => x"63000702",
          51 => x"9306f4ff",
          52 => x"63980600",
          53 => x"b387e700",
          54 => x"13041000",
          55 => x"6f000006",
          56 => x"1306f00f",
          57 => x"6318c402",
          58 => x"13f77700",
          59 => x"630a0734",
          60 => x"13f7f700",
          61 => x"93064000",
          62 => x"6304d734",
          63 => x"93874700",
          64 => x"6f000034",
          65 => x"1306f00f",
          66 => x"e300c4fe",
          67 => x"37060004",
          68 => x"3367c700",
          69 => x"9305b001",
          70 => x"13061000",
          71 => x"63ced500",
          72 => x"13060002",
          73 => x"b355d700",
          74 => x"b306d640",
          75 => x"3317d700",
          76 => x"3337e000",
          77 => x"33e6e500",
          78 => x"b387c700",
          79 => x"37070004",
          80 => x"33f7e700",
          81 => x"e30207fa",
          82 => x"13041400",
          83 => x"1307f00f",
          84 => x"6306e42e",
          85 => x"3707007e",
          86 => x"93f61700",
          87 => x"1307f7ff",
          88 => x"93d71700",
          89 => x"b3f7e700",
          90 => x"b3e7d700",
          91 => x"6ff0dff7",
          92 => x"63860606",
          93 => x"b3068540",
          94 => x"63100402",
          95 => x"6386072a",
          96 => x"1386f6ff",
          97 => x"e30806f4",
          98 => x"9305f00f",
          99 => x"6390b602",
         100 => x"93070700",
         101 => x"6f000021",
         102 => x"1306f00f",
         103 => x"e30ac5fe",
         104 => x"37060004",
         105 => x"b3e7c700",
         106 => x"13860600",
         107 => x"9305b001",
         108 => x"93061000",
         109 => x"63cec500",
         110 => x"93060002",
         111 => x"b386c640",
         112 => x"b3d5c700",
         113 => x"b397d700",
         114 => x"b337f000",
         115 => x"b3e6f500",
         116 => x"b387e600",
         117 => x"13040500",
         118 => x"6ff05ff6",
         119 => x"93061400",
         120 => x"13f6e60f",
         121 => x"63160604",
         122 => x"63180402",
         123 => x"63820724",
         124 => x"e30c07ee",
         125 => x"b387e700",
         126 => x"37070004",
         127 => x"33f7e700",
         128 => x"e30407ee",
         129 => x"370700fc",
         130 => x"1307f7ff",
         131 => x"b3f7e700",
         132 => x"13041000",
         133 => x"6ff05fed",
         134 => x"e38c07f6",
         135 => x"63040718",
         136 => x"93040000",
         137 => x"b7070002",
         138 => x"1304f00f",
         139 => x"6f004021",
         140 => x"1306f00f",
         141 => x"6382c620",
         142 => x"3387e700",
         143 => x"93571700",
         144 => x"13840600",
         145 => x"6ff05fea",
         146 => x"635ed006",
         147 => x"63120506",
         148 => x"e30c07e8",
         149 => x"9306f4ff",
         150 => x"63980600",
         151 => x"b387e740",
         152 => x"13041000",
         153 => x"6f004003",
         154 => x"1306f00f",
         155 => x"e30ec4e6",
         156 => x"9305b001",
         157 => x"13061000",
         158 => x"63ced500",
         159 => x"13060002",
         160 => x"b355d700",
         161 => x"b306d640",
         162 => x"3317d700",
         163 => x"3337e000",
         164 => x"33e6e500",
         165 => x"b387c740",
         166 => x"37090004",
         167 => x"33f72701",
         168 => x"e30407e4",
         169 => x"1309f9ff",
         170 => x"33f92701",
         171 => x"6f008011",
         172 => x"1306f00f",
         173 => x"e30ac4e2",
         174 => x"37060004",
         175 => x"3367c700",
         176 => x"6ff01ffb",
         177 => x"63800608",
         178 => x"b3068540",
         179 => x"63180402",
         180 => x"6382071e",
         181 => x"1386f6ff",
         182 => x"63180600",
         183 => x"b307f740",
         184 => x"93840500",
         185 => x"6ff0dff7",
         186 => x"1308f00f",
         187 => x"63920603",
         188 => x"93070700",
         189 => x"1304f00f",
         190 => x"6f00c006",
         191 => x"1306f00f",
         192 => x"e308c5fe",
         193 => x"37060004",
         194 => x"b3e7c700",
         195 => x"13860600",
         196 => x"1308b001",
         197 => x"93061000",
         198 => x"634ec800",
         199 => x"93060002",
         200 => x"b386c640",
         201 => x"33d8c700",
         202 => x"b397d700",
         203 => x"b337f000",
         204 => x"b366f800",
         205 => x"b307d740",
         206 => x"13040500",
         207 => x"93840500",
         208 => x"6ff09ff5",
         209 => x"93061400",
         210 => x"93f6e60f",
         211 => x"63900606",
         212 => x"63120404",
         213 => x"639c0700",
         214 => x"93040000",
         215 => x"6302070e",
         216 => x"93070700",
         217 => x"93840500",
         218 => x"6ff01fd8",
         219 => x"e30e07d6",
         220 => x"b386e740",
         221 => x"37060004",
         222 => x"33f6c600",
         223 => x"b307f740",
         224 => x"e31206fe",
         225 => x"93070000",
         226 => x"63820608",
         227 => x"93870600",
         228 => x"6ff09fd5",
         229 => x"e39407e8",
         230 => x"e30407e8",
         231 => x"93070700",
         232 => x"93840500",
         233 => x"1304f00f",
         234 => x"6ff01fd4",
         235 => x"3389e740",
         236 => x"b7060004",
         237 => x"b376d900",
         238 => x"63840604",
         239 => x"3309f740",
         240 => x"93840500",
         241 => x"13050900",
         242 => x"ef00101f",
         243 => x"1305b5ff",
         244 => x"3319a900",
         245 => x"63408504",
         246 => x"33058540",
         247 => x"13051500",
         248 => x"13070002",
         249 => x"3307a740",
         250 => x"b357a900",
         251 => x"3319e900",
         252 => x"33392001",
         253 => x"b3e72701",
         254 => x"13040000",
         255 => x"6ff0dfce",
         256 => x"e31209fc",
         257 => x"93070000",
         258 => x"13040000",
         259 => x"93040000",
         260 => x"6f000003",
         261 => x"b70700fc",
         262 => x"9387f7ff",
         263 => x"3304a440",
         264 => x"b377f900",
         265 => x"6ff05fcc",
         266 => x"93070700",
         267 => x"6ff05fe1",
         268 => x"93070700",
         269 => x"6ff05fcb",
         270 => x"1304f00f",
         271 => x"93070000",
         272 => x"37070004",
         273 => x"33f7e700",
         274 => x"630e0700",
         275 => x"13041400",
         276 => x"1307f00f",
         277 => x"6306e406",
         278 => x"370700fc",
         279 => x"1307f7ff",
         280 => x"b3f7e700",
         281 => x"1307f00f",
         282 => x"93d73700",
         283 => x"6318e400",
         284 => x"63860700",
         285 => x"b7074000",
         286 => x"93040000",
         287 => x"13147401",
         288 => x"3707807f",
         289 => x"93979700",
         290 => x"3374e400",
         291 => x"93d79700",
         292 => x"3364f400",
         293 => x"1395f401",
         294 => x"8320c100",
         295 => x"3365a400",
         296 => x"03248100",
         297 => x"83244100",
         298 => x"03290100",
         299 => x"13010101",
         300 => x"67800000",
         301 => x"93070700",
         302 => x"13840600",
         303 => x"6ff09fea",
         304 => x"93070000",
         305 => x"6ff01ffa",
         306 => x"130101fd",
         307 => x"23229102",
         308 => x"93547501",
         309 => x"232e3101",
         310 => x"232a5101",
         311 => x"23286101",
         312 => x"931a9500",
         313 => x"23261102",
         314 => x"23248102",
         315 => x"23202103",
         316 => x"232c4101",
         317 => x"23267101",
         318 => x"23248101",
         319 => x"93f4f40f",
         320 => x"138b0500",
         321 => x"93da9a00",
         322 => x"9359f501",
         323 => x"63840408",
         324 => x"9307f00f",
         325 => x"6380f40a",
         326 => x"939a3a00",
         327 => x"b7070004",
         328 => x"b3eafa00",
         329 => x"938414f8",
         330 => x"930b0000",
         331 => x"93577b01",
         332 => x"13149b00",
         333 => x"93f7f70f",
         334 => x"13549400",
         335 => x"135bfb01",
         336 => x"638a0708",
         337 => x"1307f00f",
         338 => x"6386e70a",
         339 => x"13143400",
         340 => x"37070004",
         341 => x"3364e400",
         342 => x"938717f8",
         343 => x"13070000",
         344 => x"338af440",
         345 => x"93972b00",
         346 => x"b3e7e700",
         347 => x"9387f7ff",
         348 => x"9306e000",
         349 => x"33c96901",
         350 => x"63eef608",
         351 => x"b7160000",
         352 => x"93972700",
         353 => x"9386c6f6",
         354 => x"b387d700",
         355 => x"83a70700",
         356 => x"67800700",
         357 => x"638a0a02",
         358 => x"13850a00",
         359 => x"ef00d001",
         360 => x"9307b5ff",
         361 => x"9304a0f8",
         362 => x"b39afa00",
         363 => x"b384a440",
         364 => x"6ff09ff7",
         365 => x"9304f00f",
         366 => x"930b2000",
         367 => x"e3880af6",
         368 => x"930b3000",
         369 => x"6ff09ff6",
         370 => x"93040000",
         371 => x"930b1000",
         372 => x"6ff0dff5",
         373 => x"630a0402",
         374 => x"13050400",
         375 => x"ef00c07d",
         376 => x"9307b5ff",
         377 => x"3314f400",
         378 => x"9307a0f8",
         379 => x"b387a740",
         380 => x"6ff0dff6",
         381 => x"9307f00f",
         382 => x"13072000",
         383 => x"e30204f6",
         384 => x"13073000",
         385 => x"6ff0dff5",
         386 => x"93070000",
         387 => x"13071000",
         388 => x"6ff01ff5",
         389 => x"131c5400",
         390 => x"63fa8a16",
         391 => x"130afaff",
         392 => x"13040000",
         393 => x"135b0c01",
         394 => x"b7090100",
         395 => x"93050b00",
         396 => x"9389f9ff",
         397 => x"13850a00",
         398 => x"ef00406d",
         399 => x"b3793c01",
         400 => x"93050500",
         401 => x"930b0500",
         402 => x"13850900",
         403 => x"ef004069",
         404 => x"93040500",
         405 => x"93050b00",
         406 => x"13850a00",
         407 => x"ef00806f",
         408 => x"93570401",
         409 => x"13150501",
         410 => x"b3e7a700",
         411 => x"13840b00",
         412 => x"63fe9700",
         413 => x"b3878701",
         414 => x"1384fbff",
         415 => x"63e88701",
         416 => x"63f69700",
         417 => x"1384ebff",
         418 => x"b3878701",
         419 => x"b3849740",
         420 => x"93050b00",
         421 => x"13850400",
         422 => x"ef004067",
         423 => x"93050500",
         424 => x"930a0500",
         425 => x"13850900",
         426 => x"ef008063",
         427 => x"93090500",
         428 => x"93050b00",
         429 => x"13850400",
         430 => x"ef00c069",
         431 => x"93170501",
         432 => x"13870a00",
         433 => x"63fe3701",
         434 => x"b3878701",
         435 => x"1387faff",
         436 => x"63e88701",
         437 => x"63f63701",
         438 => x"1387eaff",
         439 => x"b3878701",
         440 => x"13140401",
         441 => x"b3873741",
         442 => x"3364e400",
         443 => x"b337f000",
         444 => x"3364f400",
         445 => x"1307fa07",
         446 => x"6354e00e",
         447 => x"93777400",
         448 => x"638a0700",
         449 => x"9377f400",
         450 => x"93064000",
         451 => x"6384d700",
         452 => x"13044400",
         453 => x"b7070008",
         454 => x"b377f400",
         455 => x"638a0700",
         456 => x"b70700f8",
         457 => x"9387f7ff",
         458 => x"3374f400",
         459 => x"13070a08",
         460 => x"9307e00f",
         461 => x"63c4e708",
         462 => x"93573400",
         463 => x"8320c102",
         464 => x"03248102",
         465 => x"13177701",
         466 => x"b706807f",
         467 => x"93979700",
         468 => x"3377d700",
         469 => x"93d79700",
         470 => x"1315f901",
         471 => x"3367f700",
         472 => x"83244102",
         473 => x"03290102",
         474 => x"8329c101",
         475 => x"032a8101",
         476 => x"832a4101",
         477 => x"032b0101",
         478 => x"832bc100",
         479 => x"032c8100",
         480 => x"3365a700",
         481 => x"13010103",
         482 => x"67800000",
         483 => x"1394fa01",
         484 => x"93da1a00",
         485 => x"6ff01fe9",
         486 => x"13890900",
         487 => x"13840a00",
         488 => x"13870b00",
         489 => x"93073000",
         490 => x"6308f708",
         491 => x"93071000",
         492 => x"630cf708",
         493 => x"93072000",
         494 => x"e31ef7f2",
         495 => x"93070000",
         496 => x"1307f00f",
         497 => x"6ff09ff7",
         498 => x"13090b00",
         499 => x"6ff09ffd",
         500 => x"37044000",
         501 => x"13090000",
         502 => x"13073000",
         503 => x"6ff09ffc",
         504 => x"93071000",
         505 => x"b387e740",
         506 => x"1307b001",
         507 => x"634ef704",
         508 => x"9304ea09",
         509 => x"b357f400",
         510 => x"33149400",
         511 => x"33348000",
         512 => x"b3e78700",
         513 => x"13f77700",
         514 => x"630a0700",
         515 => x"13f7f700",
         516 => x"93064000",
         517 => x"6304d700",
         518 => x"93874700",
         519 => x"37070004",
         520 => x"33f7e700",
         521 => x"93d73700",
         522 => x"e30a07f0",
         523 => x"93070000",
         524 => x"13071000",
         525 => x"6ff09ff0",
         526 => x"b7074000",
         527 => x"1307f00f",
         528 => x"13090000",
         529 => x"6ff09fef",
         530 => x"93070000",
         531 => x"13070000",
         532 => x"6ff0dfee",
         533 => x"130101fe",
         534 => x"23282101",
         535 => x"13597501",
         536 => x"232a9100",
         537 => x"23263101",
         538 => x"23225101",
         539 => x"93149500",
         540 => x"232e1100",
         541 => x"232c8100",
         542 => x"23244101",
         543 => x"1379f90f",
         544 => x"938a0500",
         545 => x"93d49400",
         546 => x"9359f501",
         547 => x"6302091c",
         548 => x"9307f00f",
         549 => x"630ef91c",
         550 => x"93943400",
         551 => x"b7070004",
         552 => x"b3e4f400",
         553 => x"130919f8",
         554 => x"130a0000",
         555 => x"93d77a01",
         556 => x"13949a00",
         557 => x"93f7f70f",
         558 => x"13549400",
         559 => x"93dafa01",
         560 => x"6388071c",
         561 => x"1307f00f",
         562 => x"6384e71e",
         563 => x"13143400",
         564 => x"37070004",
         565 => x"3364e400",
         566 => x"938717f8",
         567 => x"93060000",
         568 => x"3309f900",
         569 => x"93172a00",
         570 => x"b3e7d700",
         571 => x"1307a000",
         572 => x"33c85901",
         573 => x"93081900",
         574 => x"6344f722",
         575 => x"13072000",
         576 => x"6348f71c",
         577 => x"9387f7ff",
         578 => x"13071000",
         579 => x"6374f71e",
         580 => x"b70e0100",
         581 => x"1383feff",
         582 => x"93df0401",
         583 => x"135f0401",
         584 => x"b3f46400",
         585 => x"33746400",
         586 => x"13850400",
         587 => x"93050400",
         588 => x"ef00003b",
         589 => x"13070500",
         590 => x"93050f00",
         591 => x"13850400",
         592 => x"ef00003a",
         593 => x"93070500",
         594 => x"93050400",
         595 => x"13850f00",
         596 => x"ef000039",
         597 => x"130e0500",
         598 => x"93050f00",
         599 => x"13850f00",
         600 => x"ef000038",
         601 => x"13540701",
         602 => x"b387c701",
         603 => x"3304f400",
         604 => x"93060500",
         605 => x"6374c401",
         606 => x"b306d501",
         607 => x"b3776400",
         608 => x"33776700",
         609 => x"93970701",
         610 => x"b387e700",
         611 => x"13976700",
         612 => x"13540401",
         613 => x"3337e000",
         614 => x"93d7a701",
         615 => x"3304d400",
         616 => x"b367f700",
         617 => x"13146400",
         618 => x"3364f400",
         619 => x"b7070008",
         620 => x"b377f400",
         621 => x"638e0718",
         622 => x"93571400",
         623 => x"13741400",
         624 => x"33e48700",
         625 => x"1387f807",
         626 => x"6358e018",
         627 => x"93777400",
         628 => x"638a0700",
         629 => x"9377f400",
         630 => x"93064000",
         631 => x"6384d700",
         632 => x"13044400",
         633 => x"b7070008",
         634 => x"b377f400",
         635 => x"638a0700",
         636 => x"b70700f8",
         637 => x"9387f7ff",
         638 => x"3374f400",
         639 => x"13870808",
         640 => x"9307e00f",
         641 => x"63cee71a",
         642 => x"93573400",
         643 => x"8320c101",
         644 => x"03248101",
         645 => x"13177701",
         646 => x"b706807f",
         647 => x"93979700",
         648 => x"3377d700",
         649 => x"93d79700",
         650 => x"3367f700",
         651 => x"1315f801",
         652 => x"83244101",
         653 => x"03290101",
         654 => x"8329c100",
         655 => x"032a8100",
         656 => x"832a4100",
         657 => x"3365a700",
         658 => x"13010102",
         659 => x"67800000",
         660 => x"638a0402",
         661 => x"13850400",
         662 => x"ef000036",
         663 => x"9307b5ff",
         664 => x"1309a0f8",
         665 => x"b394f400",
         666 => x"3309a940",
         667 => x"6ff0dfe3",
         668 => x"1309f00f",
         669 => x"130a2000",
         670 => x"e38a04e2",
         671 => x"130a3000",
         672 => x"6ff0dfe2",
         673 => x"13090000",
         674 => x"130a1000",
         675 => x"6ff01fe2",
         676 => x"630a0402",
         677 => x"13050400",
         678 => x"ef000032",
         679 => x"9307b5ff",
         680 => x"3314f400",
         681 => x"9307a0f8",
         682 => x"b387a740",
         683 => x"6ff01fe3",
         684 => x"9307f00f",
         685 => x"93062000",
         686 => x"e30404e2",
         687 => x"93063000",
         688 => x"6ff01fe2",
         689 => x"93070000",
         690 => x"93061000",
         691 => x"6ff05fe1",
         692 => x"13071000",
         693 => x"b317f700",
         694 => x"13f70753",
         695 => x"631c0704",
         696 => x"13f70724",
         697 => x"6316070c",
         698 => x"93f78708",
         699 => x"e38207e2",
         700 => x"13880a00",
         701 => x"13062000",
         702 => x"93070000",
         703 => x"1307f00f",
         704 => x"e386c6f0",
         705 => x"93073000",
         706 => x"6384f60a",
         707 => x"93071000",
         708 => x"e39af6ea",
         709 => x"93070000",
         710 => x"13070000",
         711 => x"6ff01fef",
         712 => x"1307f000",
         713 => x"638ee700",
         714 => x"1307b000",
         715 => x"e382e7fc",
         716 => x"13880900",
         717 => x"13840400",
         718 => x"93060a00",
         719 => x"6ff09ffb",
         720 => x"37044000",
         721 => x"13080000",
         722 => x"93063000",
         723 => x"6ff09ffb",
         724 => x"93080900",
         725 => x"6ff01fe7",
         726 => x"93071000",
         727 => x"b387e740",
         728 => x"1307b001",
         729 => x"e348f7fa",
         730 => x"9388e809",
         731 => x"b357f400",
         732 => x"33141401",
         733 => x"33348000",
         734 => x"b3e78700",
         735 => x"13f77700",
         736 => x"630a0700",
         737 => x"13f7f700",
         738 => x"93064000",
         739 => x"6304d700",
         740 => x"93874700",
         741 => x"37070004",
         742 => x"33f7e700",
         743 => x"93d73700",
         744 => x"e30607e6",
         745 => x"93070000",
         746 => x"13071000",
         747 => x"6ff01fe6",
         748 => x"b7074000",
         749 => x"1307f00f",
         750 => x"13080000",
         751 => x"6ff01fe5",
         752 => x"93070000",
         753 => x"1307f00f",
         754 => x"6ff05fe4",
         755 => x"6308050e",
         756 => x"9357f541",
         757 => x"130101ff",
         758 => x"23248100",
         759 => x"33c4a700",
         760 => x"3304f440",
         761 => x"23229100",
         762 => x"9354f501",
         763 => x"13050400",
         764 => x"23261100",
         765 => x"ef00401c",
         766 => x"1307e009",
         767 => x"3307a740",
         768 => x"93076009",
         769 => x"63cce702",
         770 => x"130585ff",
         771 => x"b317a400",
         772 => x"8320c100",
         773 => x"03248100",
         774 => x"93979700",
         775 => x"13177701",
         776 => x"93d79700",
         777 => x"1395f401",
         778 => x"3367f700",
         779 => x"83244100",
         780 => x"3365a700",
         781 => x"13010101",
         782 => x"67800000",
         783 => x"93079009",
         784 => x"63d0e702",
         785 => x"93075000",
         786 => x"b387a740",
         787 => x"9306b501",
         788 => x"b357f400",
         789 => x"3314d400",
         790 => x"33348000",
         791 => x"33e48700",
         792 => x"93075000",
         793 => x"63d6a700",
         794 => x"9307b5ff",
         795 => x"3314f400",
         796 => x"b70700fc",
         797 => x"9387f7ff",
         798 => x"93767400",
         799 => x"b377f400",
         800 => x"638a0600",
         801 => x"1374f400",
         802 => x"93064000",
         803 => x"6304d400",
         804 => x"93874700",
         805 => x"b7060004",
         806 => x"b3f6d700",
         807 => x"638c0600",
         808 => x"370700fc",
         809 => x"1307f7ff",
         810 => x"b3f7e700",
         811 => x"1307f009",
         812 => x"3307a740",
         813 => x"93d73700",
         814 => x"6ff09ff5",
         815 => x"93070000",
         816 => x"13070000",
         817 => x"93979700",
         818 => x"93d79700",
         819 => x"13177701",
         820 => x"3367f700",
         821 => x"1315f501",
         822 => x"3365a700",
         823 => x"67800000",
         824 => x"13060500",
         825 => x"13050000",
         826 => x"93f61500",
         827 => x"63840600",
         828 => x"3305c500",
         829 => x"93d51500",
         830 => x"13161600",
         831 => x"e39605fe",
         832 => x"67800000",
         833 => x"63400506",
         834 => x"63c60506",
         835 => x"13860500",
         836 => x"93050500",
         837 => x"1305f0ff",
         838 => x"630c0602",
         839 => x"93061000",
         840 => x"637ab600",
         841 => x"6358c000",
         842 => x"13161600",
         843 => x"93961600",
         844 => x"e36ab6fe",
         845 => x"13050000",
         846 => x"63e6c500",
         847 => x"b385c540",
         848 => x"3365d500",
         849 => x"93d61600",
         850 => x"13561600",
         851 => x"e39606fe",
         852 => x"67800000",
         853 => x"93820000",
         854 => x"eff05ffb",
         855 => x"13850500",
         856 => x"67800200",
         857 => x"3305a040",
         858 => x"6348b000",
         859 => x"b305b040",
         860 => x"6ff0dff9",
         861 => x"b305b040",
         862 => x"93820000",
         863 => x"eff01ff9",
         864 => x"3305a040",
         865 => x"67800200",
         866 => x"93820000",
         867 => x"63ca0500",
         868 => x"634c0500",
         869 => x"eff09ff7",
         870 => x"13850500",
         871 => x"67800200",
         872 => x"b305b040",
         873 => x"e35805fe",
         874 => x"3305a040",
         875 => x"eff01ff6",
         876 => x"3305b040",
         877 => x"67800200",
         878 => x"b7070100",
         879 => x"637af502",
         880 => x"93370510",
         881 => x"93c71700",
         882 => x"93973700",
         883 => x"37170000",
         884 => x"93060002",
         885 => x"b386f640",
         886 => x"3355f500",
         887 => x"930787fa",
         888 => x"b387a700",
         889 => x"03c50700",
         890 => x"3385a640",
         891 => x"67800000",
         892 => x"37070001",
         893 => x"93070001",
         894 => x"e36ae5fc",
         895 => x"93078001",
         896 => x"6ff0dffc",
         897 => x"130101fe",
         898 => x"b7170000",
         899 => x"23225101",
         900 => x"83aa870a",
         901 => x"232c8100",
         902 => x"232a9100",
         903 => x"23282101",
         904 => x"23244101",
         905 => x"232e1100",
         906 => x"23263101",
         907 => x"13041000",
         908 => x"130a4001",
         909 => x"83a50186",
         910 => x"83a94186",
         911 => x"13850a00",
         912 => x"eff08fe8",
         913 => x"93850900",
         914 => x"eff0cfa2",
         915 => x"23a2a186",
         916 => x"83a90186",
         917 => x"13050400",
         918 => x"eff05fd7",
         919 => x"93850900",
         920 => x"eff05f9f",
         921 => x"13041400",
         922 => x"23a0a186",
         923 => x"e31444fd",
         924 => x"8320c101",
         925 => x"03248101",
         926 => x"83244101",
         927 => x"03290101",
         928 => x"8329c100",
         929 => x"032a8100",
         930 => x"832a4100",
         931 => x"13050000",
         932 => x"13010102",
         933 => x"67800000",
         934 => x"130101ff",
         935 => x"23248100",
         936 => x"23229100",
         937 => x"37140000",
         938 => x"b7140000",
         939 => x"9387040b",
         940 => x"1304040b",
         941 => x"3304f440",
         942 => x"23202101",
         943 => x"23261100",
         944 => x"13542440",
         945 => x"9384040b",
         946 => x"13090000",
         947 => x"63108904",
         948 => x"b7140000",
         949 => x"37140000",
         950 => x"9387040b",
         951 => x"1304040b",
         952 => x"3304f440",
         953 => x"13542440",
         954 => x"9384040b",
         955 => x"13090000",
         956 => x"63188902",
         957 => x"8320c100",
         958 => x"03248100",
         959 => x"83244100",
         960 => x"03290100",
         961 => x"13010101",
         962 => x"67800000",
         963 => x"83a70400",
         964 => x"13091900",
         965 => x"93844400",
         966 => x"e7800700",
         967 => x"6ff01ffb",
         968 => x"83a70400",
         969 => x"13091900",
         970 => x"93844400",
         971 => x"e7800700",
         972 => x"6ff01ffc",
         973 => x"9308d005",
         974 => x"73000000",
         975 => x"63520502",
         976 => x"130101ff",
         977 => x"23248100",
         978 => x"13040500",
         979 => x"23261100",
         980 => x"33048040",
         981 => x"ef000001",
         982 => x"23208500",
         983 => x"6f000000",
         984 => x"6f000000",
         985 => x"03a58186",
         986 => x"67800000",
         987 => x"bc070000",
         988 => x"48080000",
         989 => x"c8070000",
         990 => x"48080000",
         991 => x"38080000",
         992 => x"48080000",
         993 => x"c8070000",
         994 => x"bc070000",
         995 => x"bc070000",
         996 => x"38080000",
         997 => x"c8070000",
         998 => x"98070000",
         999 => x"98070000",
        1000 => x"98070000",
        1001 => x"d0070000",
        1002 => x"00010202",
        1003 => x"03030303",
        1004 => x"04040404",
        1005 => x"04040404",
        1006 => x"05050505",
        1007 => x"05050505",
        1008 => x"05050505",
        1009 => x"05050505",
        1010 => x"06060606",
        1011 => x"06060606",
        1012 => x"06060606",
        1013 => x"06060606",
        1014 => x"06060606",
        1015 => x"06060606",
        1016 => x"06060606",
        1017 => x"06060606",
        1018 => x"07070707",
        1019 => x"07070707",
        1020 => x"07070707",
        1021 => x"07070707",
        1022 => x"07070707",
        1023 => x"07070707",
        1024 => x"07070707",
        1025 => x"07070707",
        1026 => x"07070707",
        1027 => x"07070707",
        1028 => x"07070707",
        1029 => x"07070707",
        1030 => x"07070707",
        1031 => x"07070707",
        1032 => x"07070707",
        1033 => x"07070707",
        1034 => x"08080808",
        1035 => x"08080808",
        1036 => x"08080808",
        1037 => x"08080808",
        1038 => x"08080808",
        1039 => x"08080808",
        1040 => x"08080808",
        1041 => x"08080808",
        1042 => x"08080808",
        1043 => x"08080808",
        1044 => x"08080808",
        1045 => x"08080808",
        1046 => x"08080808",
        1047 => x"08080808",
        1048 => x"08080808",
        1049 => x"08080808",
        1050 => x"08080808",
        1051 => x"08080808",
        1052 => x"08080808",
        1053 => x"08080808",
        1054 => x"08080808",
        1055 => x"08080808",
        1056 => x"08080808",
        1057 => x"08080808",
        1058 => x"08080808",
        1059 => x"08080808",
        1060 => x"08080808",
        1061 => x"08080808",
        1062 => x"08080808",
        1063 => x"08080808",
        1064 => x"08080808",
        1065 => x"08080808",
        1066 => x"0000803f",
        1067 => x"00000020",
        1068 => x"00000000",
        1069 => x"00000000",
        1070 => x"00000000",
        1071 => x"00000000",
        1072 => x"00000000",
        1073 => x"00000000",
        1074 => x"00000000",
        1075 => x"00000000",
        1076 => x"00000000",
        1077 => x"00000000",
        1078 => x"00000000",
        1079 => x"00000000",
        1080 => x"00000000",
        1081 => x"00000000",
        1082 => x"00000000",
        1083 => x"00000000",
        1084 => x"00000000",
        1085 => x"00000000",
        1086 => x"00000000",
        1087 => x"00000000",
        1088 => x"00000000",
        1089 => x"00000000",
        1090 => x"00000000",
        1091 => x"00000000",
        1092 => x"0000803f",
        1093 => x"0000803f",
        1094 => x"00000020",
        others => (others => '0')
    );
end package processor_common_rom;
