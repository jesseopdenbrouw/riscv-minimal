-- srec2vhdl table generator
-- for input file main.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"93828206",
           6 => x"73905230",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef10803c",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"938585fd",
          21 => x"13050500",
          22 => x"ef100038",
          23 => x"ef10406f",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10403e",
          29 => x"ef10c069",
          30 => x"6f000000",
          31 => x"37170000",
          32 => x"b70700f0",
          33 => x"13077745",
          34 => x"23a2e702",
          35 => x"13070004",
          36 => x"23a4e702",
          37 => x"67800000",
          38 => x"1375f50f",
          39 => x"b70700f0",
          40 => x"23a0a702",
          41 => x"370700f0",
          42 => x"8327c702",
          43 => x"93f70701",
          44 => x"e38c07fe",
          45 => x"67800000",
          46 => x"63060502",
          47 => x"83470500",
          48 => x"63820702",
          49 => x"370700f0",
          50 => x"13051500",
          51 => x"2320f702",
          52 => x"8327c702",
          53 => x"93f70701",
          54 => x"e38c07fe",
          55 => x"83470500",
          56 => x"e39407fe",
          57 => x"67800000",
          58 => x"370700f0",
          59 => x"8327c702",
          60 => x"93f74700",
          61 => x"e38c07fe",
          62 => x"03250702",
          63 => x"1375f50f",
          64 => x"67800000",
          65 => x"130101ff",
          66 => x"373e0000",
          67 => x"370700f0",
          68 => x"930e0500",
          69 => x"138ff5ff",
          70 => x"23268100",
          71 => x"13050000",
          72 => x"130ecebd",
          73 => x"13070702",
          74 => x"13035001",
          75 => x"93027000",
          76 => x"930fe005",
          77 => x"9305f007",
          78 => x"93082000",
          79 => x"13082001",
          80 => x"b7330000",
          81 => x"1306f007",
          82 => x"8327c700",
          83 => x"93f74700",
          84 => x"e38c07fe",
          85 => x"03240700",
          86 => x"9376f40f",
          87 => x"636ed302",
          88 => x"63fed802",
          89 => x"9387d6ff",
          90 => x"636af802",
          91 => x"93972700",
          92 => x"b307fe00",
          93 => x"83a70700",
          94 => x"67800700",
          95 => x"1305f5ff",
          96 => x"6308050c",
          97 => x"2320c700",
          98 => x"8327c700",
          99 => x"93f70701",
         100 => x"e38c07fe",
         101 => x"6ff09ffe",
         102 => x"638cb606",
         103 => x"635ae50d",
         104 => x"1374f40f",
         105 => x"930704fe",
         106 => x"93f7f70f",
         107 => x"e3eefff8",
         108 => x"b387ae00",
         109 => x"23808700",
         110 => x"13051500",
         111 => x"2320d700",
         112 => x"8327c700",
         113 => x"93f70701",
         114 => x"e38c07fe",
         115 => x"6ff0dff7",
         116 => x"b38eae00",
         117 => x"b7360000",
         118 => x"23800e00",
         119 => x"9307d000",
         120 => x"938686e5",
         121 => x"370700f0",
         122 => x"93861600",
         123 => x"2320f702",
         124 => x"8327c702",
         125 => x"93f70701",
         126 => x"e38c07fe",
         127 => x"83c70600",
         128 => x"e39407fe",
         129 => x"0324c100",
         130 => x"13010101",
         131 => x"67800000",
         132 => x"63040504",
         133 => x"2320b700",
         134 => x"8327c700",
         135 => x"93f70701",
         136 => x"e38c07fe",
         137 => x"1305f5ff",
         138 => x"6ff01ff2",
         139 => x"9307c003",
         140 => x"938603f2",
         141 => x"93861600",
         142 => x"2320f700",
         143 => x"8327c700",
         144 => x"93f70701",
         145 => x"e38c07fe",
         146 => x"83c70600",
         147 => x"e39407fe",
         148 => x"13050000",
         149 => x"6ff05fef",
         150 => x"23205700",
         151 => x"8327c700",
         152 => x"93f70701",
         153 => x"e38c07fe",
         154 => x"13050000",
         155 => x"6ff0dfed",
         156 => x"23205700",
         157 => x"8327c700",
         158 => x"93f70701",
         159 => x"e38c07fe",
         160 => x"6ff09fec",
         161 => x"1375f50f",
         162 => x"b70700f0",
         163 => x"23a0a702",
         164 => x"370700f0",
         165 => x"8327c702",
         166 => x"93f70701",
         167 => x"e38c07fe",
         168 => x"13051000",
         169 => x"67800000",
         170 => x"370700f0",
         171 => x"8327c702",
         172 => x"93f74700",
         173 => x"e38c07fe",
         174 => x"03250702",
         175 => x"1375f50f",
         176 => x"67800000",
         177 => x"13050000",
         178 => x"67800000",
         179 => x"13050000",
         180 => x"67800000",
         181 => x"130101f8",
         182 => x"23221100",
         183 => x"23242100",
         184 => x"23263100",
         185 => x"23284100",
         186 => x"232a5100",
         187 => x"232c6100",
         188 => x"232e7100",
         189 => x"23208102",
         190 => x"23229102",
         191 => x"2324a102",
         192 => x"2326b102",
         193 => x"2328c102",
         194 => x"232ad102",
         195 => x"232ce102",
         196 => x"232ef102",
         197 => x"23200105",
         198 => x"23221105",
         199 => x"23242105",
         200 => x"23263105",
         201 => x"23284105",
         202 => x"232a5105",
         203 => x"232c6105",
         204 => x"232e7105",
         205 => x"23208107",
         206 => x"23229107",
         207 => x"2324a107",
         208 => x"2326b107",
         209 => x"2328c107",
         210 => x"232ad107",
         211 => x"232ce107",
         212 => x"232ef107",
         213 => x"f3272034",
         214 => x"37070080",
         215 => x"93067700",
         216 => x"6388d70c",
         217 => x"9306b000",
         218 => x"63e4f602",
         219 => x"13071000",
         220 => x"637cf70a",
         221 => x"63eaf60a",
         222 => x"37370000",
         223 => x"93972700",
         224 => x"130787c2",
         225 => x"b387e700",
         226 => x"83a70700",
         227 => x"67800700",
         228 => x"93061701",
         229 => x"6384d70a",
         230 => x"13072701",
         231 => x"6396e708",
         232 => x"ef008038",
         233 => x"03258102",
         234 => x"832fc107",
         235 => x"032f8107",
         236 => x"832e4107",
         237 => x"032e0107",
         238 => x"832dc106",
         239 => x"032d8106",
         240 => x"832c4106",
         241 => x"032c0106",
         242 => x"832bc105",
         243 => x"032b8105",
         244 => x"832a4105",
         245 => x"032a0105",
         246 => x"8329c104",
         247 => x"03298104",
         248 => x"83284104",
         249 => x"03280104",
         250 => x"8327c103",
         251 => x"03278103",
         252 => x"83264103",
         253 => x"03260103",
         254 => x"8325c102",
         255 => x"83244102",
         256 => x"03240102",
         257 => x"8323c101",
         258 => x"03238101",
         259 => x"83224101",
         260 => x"03220101",
         261 => x"8321c100",
         262 => x"03218100",
         263 => x"83204100",
         264 => x"13010108",
         265 => x"73002030",
         266 => x"03258102",
         267 => x"6ff0dff7",
         268 => x"ef00c02a",
         269 => x"03258102",
         270 => x"6ff01ff7",
         271 => x"ef00c026",
         272 => x"03258102",
         273 => x"6ff05ff6",
         274 => x"9307600d",
         275 => x"6388f814",
         276 => x"9307900a",
         277 => x"6382f818",
         278 => x"63cc1703",
         279 => x"938878fc",
         280 => x"93074002",
         281 => x"63e81705",
         282 => x"b7370000",
         283 => x"938787c5",
         284 => x"93982800",
         285 => x"b388f800",
         286 => x"83a70800",
         287 => x"67800700",
         288 => x"13050100",
         289 => x"ef00c01b",
         290 => x"03258102",
         291 => x"6ff0dff1",
         292 => x"938808c0",
         293 => x"9307f000",
         294 => x"63ee1701",
         295 => x"b7370000",
         296 => x"9387c7ce",
         297 => x"93982800",
         298 => x"b388f800",
         299 => x"83a70800",
         300 => x"67800700",
         301 => x"ef104025",
         302 => x"93078005",
         303 => x"2320f500",
         304 => x"9307f0ff",
         305 => x"13850700",
         306 => x"6ff01fee",
         307 => x"b7270000",
         308 => x"23a2f500",
         309 => x"93070000",
         310 => x"13850700",
         311 => x"6ff0dfec",
         312 => x"93070000",
         313 => x"13850700",
         314 => x"6ff01fec",
         315 => x"ef10c021",
         316 => x"93079000",
         317 => x"2320f500",
         318 => x"9307f0ff",
         319 => x"13850700",
         320 => x"6ff09fea",
         321 => x"ef104020",
         322 => x"9307f001",
         323 => x"2320f500",
         324 => x"9307f0ff",
         325 => x"13850700",
         326 => x"6ff01fe9",
         327 => x"ef10c01e",
         328 => x"9307d000",
         329 => x"2320f500",
         330 => x"9307f0ff",
         331 => x"13850700",
         332 => x"6ff09fe7",
         333 => x"ef10401d",
         334 => x"93072000",
         335 => x"2320f500",
         336 => x"9307f0ff",
         337 => x"13850700",
         338 => x"6ff01fe6",
         339 => x"13090600",
         340 => x"13840500",
         341 => x"635cc000",
         342 => x"b384c500",
         343 => x"03450400",
         344 => x"13041400",
         345 => x"eff01fd2",
         346 => x"e39a84fe",
         347 => x"13050900",
         348 => x"6ff09fe3",
         349 => x"13090600",
         350 => x"13840500",
         351 => x"e358c0fe",
         352 => x"b384c500",
         353 => x"eff05fd2",
         354 => x"2300a400",
         355 => x"13041400",
         356 => x"e31a94fe",
         357 => x"13050900",
         358 => x"6ff01fe1",
         359 => x"63180500",
         360 => x"13858189",
         361 => x"13050500",
         362 => x"6ff01fe0",
         363 => x"b7870020",
         364 => x"93870700",
         365 => x"13070040",
         366 => x"b387e740",
         367 => x"e364f5fe",
         368 => x"ef108014",
         369 => x"9307c000",
         370 => x"2320f500",
         371 => x"1305f0ff",
         372 => x"13050500",
         373 => x"6ff05fdd",
         374 => x"13090000",
         375 => x"93040500",
         376 => x"13040900",
         377 => x"93090900",
         378 => x"93070900",
         379 => x"732410c8",
         380 => x"f32910c0",
         381 => x"f32710c8",
         382 => x"e31af4fe",
         383 => x"37460f00",
         384 => x"13060624",
         385 => x"93060000",
         386 => x"13850900",
         387 => x"93050400",
         388 => x"ef00501e",
         389 => x"37460f00",
         390 => x"23a4a400",
         391 => x"13060624",
         392 => x"93060000",
         393 => x"13850900",
         394 => x"93050400",
         395 => x"ef008059",
         396 => x"23a0a400",
         397 => x"23a2b400",
         398 => x"13050900",
         399 => x"6ff0dfd6",
         400 => x"37350000",
         401 => x"130101ff",
         402 => x"1305c5f2",
         403 => x"23261100",
         404 => x"23248100",
         405 => x"23229100",
         406 => x"23202101",
         407 => x"eff0dfa5",
         408 => x"73294034",
         409 => x"93040002",
         410 => x"37040080",
         411 => x"33758900",
         412 => x"3335a000",
         413 => x"13050503",
         414 => x"9384f4ff",
         415 => x"eff0dfa1",
         416 => x"13541400",
         417 => x"e39404fe",
         418 => x"03248100",
         419 => x"8320c100",
         420 => x"83244100",
         421 => x"03290100",
         422 => x"37350000",
         423 => x"130585e5",
         424 => x"13010101",
         425 => x"6ff05fa1",
         426 => x"b70700f0",
         427 => x"03a74708",
         428 => x"1377f7fe",
         429 => x"23a2e708",
         430 => x"03a74700",
         431 => x"13471700",
         432 => x"23a2e700",
         433 => x"67800000",
         434 => x"370700f0",
         435 => x"83274700",
         436 => x"93e70720",
         437 => x"2322f700",
         438 => x"6f000000",
         439 => x"b70700f0",
         440 => x"83a6470f",
         441 => x"03a6070f",
         442 => x"03a7470f",
         443 => x"e31ad7fe",
         444 => x"b7860100",
         445 => x"9305f0ff",
         446 => x"9386066a",
         447 => x"23aeb70e",
         448 => x"b306d600",
         449 => x"23acb70e",
         450 => x"33b6c600",
         451 => x"23acd70e",
         452 => x"3306e600",
         453 => x"23aec70e",
         454 => x"03a74700",
         455 => x"13472700",
         456 => x"23a2e700",
         457 => x"67800000",
         458 => x"370700f0",
         459 => x"8327c702",
         460 => x"93f74700",
         461 => x"638a0700",
         462 => x"83274700",
         463 => x"93c74700",
         464 => x"2322f700",
         465 => x"83270702",
         466 => x"67800000",
         467 => x"13030500",
         468 => x"138e0500",
         469 => x"93080000",
         470 => x"63dc0500",
         471 => x"b337a000",
         472 => x"330eb040",
         473 => x"330efe40",
         474 => x"3303a040",
         475 => x"9308f0ff",
         476 => x"63dc0600",
         477 => x"b337c000",
         478 => x"b306d040",
         479 => x"93c8f8ff",
         480 => x"b386f640",
         481 => x"3306c040",
         482 => x"13070600",
         483 => x"13080300",
         484 => x"93070e00",
         485 => x"639c0628",
         486 => x"b7350000",
         487 => x"9385c5d2",
         488 => x"6376ce0e",
         489 => x"b7060100",
         490 => x"6378d60c",
         491 => x"93360610",
         492 => x"93c61600",
         493 => x"93963600",
         494 => x"3355d600",
         495 => x"b385a500",
         496 => x"83c50500",
         497 => x"13050002",
         498 => x"b386d500",
         499 => x"b305d540",
         500 => x"630cd500",
         501 => x"b317be00",
         502 => x"b356d300",
         503 => x"3317b600",
         504 => x"b3e7f600",
         505 => x"3318b300",
         506 => x"93550701",
         507 => x"33deb702",
         508 => x"13160701",
         509 => x"13560601",
         510 => x"b3f7b702",
         511 => x"13050e00",
         512 => x"3303c603",
         513 => x"93960701",
         514 => x"93570801",
         515 => x"b3e7d700",
         516 => x"63fe6700",
         517 => x"b387e700",
         518 => x"1305feff",
         519 => x"63e8e700",
         520 => x"63f66700",
         521 => x"1305eeff",
         522 => x"b387e700",
         523 => x"b3876740",
         524 => x"33d3b702",
         525 => x"13180801",
         526 => x"13580801",
         527 => x"b3f7b702",
         528 => x"b3066602",
         529 => x"93970701",
         530 => x"3368f800",
         531 => x"93070300",
         532 => x"637cd800",
         533 => x"33080701",
         534 => x"9307f3ff",
         535 => x"6366e800",
         536 => x"6374d800",
         537 => x"9307e3ff",
         538 => x"13150501",
         539 => x"3365f500",
         540 => x"93050000",
         541 => x"6f00000e",
         542 => x"37050001",
         543 => x"93060001",
         544 => x"e36ca6f2",
         545 => x"93068001",
         546 => x"6ff01ff3",
         547 => x"63140600",
         548 => x"73001000",
         549 => x"b7070100",
         550 => x"637af60c",
         551 => x"93360610",
         552 => x"93c61600",
         553 => x"93963600",
         554 => x"b357d600",
         555 => x"b385f500",
         556 => x"83c70500",
         557 => x"b387d700",
         558 => x"93060002",
         559 => x"b385f640",
         560 => x"6390f60c",
         561 => x"b307ce40",
         562 => x"93051000",
         563 => x"13530701",
         564 => x"b3de6702",
         565 => x"13160701",
         566 => x"13560601",
         567 => x"93560801",
         568 => x"b3f76702",
         569 => x"13850e00",
         570 => x"330ed603",
         571 => x"93970701",
         572 => x"b3e7f600",
         573 => x"63fec701",
         574 => x"b387e700",
         575 => x"1385feff",
         576 => x"63e8e700",
         577 => x"63f6c701",
         578 => x"1385eeff",
         579 => x"b387e700",
         580 => x"b387c741",
         581 => x"33de6702",
         582 => x"13180801",
         583 => x"13580801",
         584 => x"b3f76702",
         585 => x"b306c603",
         586 => x"93970701",
         587 => x"3368f800",
         588 => x"93070e00",
         589 => x"637cd800",
         590 => x"33080701",
         591 => x"9307feff",
         592 => x"6366e800",
         593 => x"6374d800",
         594 => x"9307eeff",
         595 => x"13150501",
         596 => x"3365f500",
         597 => x"638a0800",
         598 => x"b337a000",
         599 => x"b305b040",
         600 => x"b385f540",
         601 => x"3305a040",
         602 => x"67800000",
         603 => x"b7070001",
         604 => x"93060001",
         605 => x"e36af6f2",
         606 => x"93068001",
         607 => x"6ff0dff2",
         608 => x"3317b600",
         609 => x"b356fe00",
         610 => x"13550701",
         611 => x"331ebe00",
         612 => x"b357f300",
         613 => x"b3e7c701",
         614 => x"33dea602",
         615 => x"13160701",
         616 => x"13560601",
         617 => x"3318b300",
         618 => x"b3f6a602",
         619 => x"3303c603",
         620 => x"93950601",
         621 => x"93d60701",
         622 => x"b3e6b600",
         623 => x"93050e00",
         624 => x"63fe6600",
         625 => x"b386e600",
         626 => x"9305feff",
         627 => x"63e8e600",
         628 => x"63f66600",
         629 => x"9305eeff",
         630 => x"b386e600",
         631 => x"b3866640",
         632 => x"33d3a602",
         633 => x"93970701",
         634 => x"93d70701",
         635 => x"b3f6a602",
         636 => x"33066602",
         637 => x"93960601",
         638 => x"b3e7d700",
         639 => x"93060300",
         640 => x"63fec700",
         641 => x"b387e700",
         642 => x"9306f3ff",
         643 => x"63e8e700",
         644 => x"63f6c700",
         645 => x"9306e3ff",
         646 => x"b387e700",
         647 => x"93950501",
         648 => x"b387c740",
         649 => x"b3e5d500",
         650 => x"6ff05fea",
         651 => x"6366de18",
         652 => x"b7070100",
         653 => x"63f4f604",
         654 => x"13b70610",
         655 => x"13471700",
         656 => x"13173700",
         657 => x"b7370000",
         658 => x"b3d5e600",
         659 => x"9387c7d2",
         660 => x"b387b700",
         661 => x"83c70700",
         662 => x"b387e700",
         663 => x"13070002",
         664 => x"b305f740",
         665 => x"6316f702",
         666 => x"13051000",
         667 => x"e3e4c6ef",
         668 => x"3335c300",
         669 => x"13451500",
         670 => x"6ff0dfed",
         671 => x"b7070001",
         672 => x"13070001",
         673 => x"e3e0f6fc",
         674 => x"13078001",
         675 => x"6ff09ffb",
         676 => x"3357f600",
         677 => x"b396b600",
         678 => x"b366d700",
         679 => x"3357fe00",
         680 => x"331ebe00",
         681 => x"b357f300",
         682 => x"b3e7c701",
         683 => x"13de0601",
         684 => x"335fc703",
         685 => x"13980601",
         686 => x"13580801",
         687 => x"3316b600",
         688 => x"3377c703",
         689 => x"b30ee803",
         690 => x"13150701",
         691 => x"13d70701",
         692 => x"3367a700",
         693 => x"13050f00",
         694 => x"637ed701",
         695 => x"3307d700",
         696 => x"1305ffff",
         697 => x"6368d700",
         698 => x"6376d701",
         699 => x"1305efff",
         700 => x"3307d700",
         701 => x"3307d741",
         702 => x"b35ec703",
         703 => x"93970701",
         704 => x"93d70701",
         705 => x"3377c703",
         706 => x"3308d803",
         707 => x"13170701",
         708 => x"b3e7e700",
         709 => x"13870e00",
         710 => x"63fe0701",
         711 => x"b387d700",
         712 => x"1387feff",
         713 => x"63e8d700",
         714 => x"63f60701",
         715 => x"1387eeff",
         716 => x"b387d700",
         717 => x"13150501",
         718 => x"b70e0100",
         719 => x"3365e500",
         720 => x"9386feff",
         721 => x"3377d500",
         722 => x"b3870741",
         723 => x"b376d600",
         724 => x"13580501",
         725 => x"13560601",
         726 => x"330ed702",
         727 => x"b306d802",
         728 => x"3307c702",
         729 => x"3308c802",
         730 => x"3306d700",
         731 => x"13570e01",
         732 => x"3307c700",
         733 => x"6374d700",
         734 => x"3308d801",
         735 => x"93560701",
         736 => x"b3860601",
         737 => x"63e6d702",
         738 => x"e394d7ce",
         739 => x"b7070100",
         740 => x"9387f7ff",
         741 => x"3377f700",
         742 => x"13170701",
         743 => x"337efe00",
         744 => x"3313b300",
         745 => x"3307c701",
         746 => x"93050000",
         747 => x"e374e3da",
         748 => x"1305f5ff",
         749 => x"6ff0dfcb",
         750 => x"93050000",
         751 => x"13050000",
         752 => x"6ff05fd9",
         753 => x"13030500",
         754 => x"93880500",
         755 => x"13070600",
         756 => x"13080500",
         757 => x"93870500",
         758 => x"63920628",
         759 => x"b7350000",
         760 => x"9385c5d2",
         761 => x"63f6c80e",
         762 => x"b7060100",
         763 => x"6378d60c",
         764 => x"93360610",
         765 => x"93c61600",
         766 => x"93963600",
         767 => x"3355d600",
         768 => x"b385a500",
         769 => x"83c50500",
         770 => x"13050002",
         771 => x"b386d500",
         772 => x"b305d540",
         773 => x"630cd500",
         774 => x"b397b800",
         775 => x"b356d300",
         776 => x"3317b600",
         777 => x"b3e7f600",
         778 => x"3318b300",
         779 => x"93550701",
         780 => x"33d3b702",
         781 => x"13160701",
         782 => x"13560601",
         783 => x"b3f7b702",
         784 => x"13050300",
         785 => x"b3086602",
         786 => x"93960701",
         787 => x"93570801",
         788 => x"b3e7d700",
         789 => x"63fe1701",
         790 => x"b387e700",
         791 => x"1305f3ff",
         792 => x"63e8e700",
         793 => x"63f61701",
         794 => x"1305e3ff",
         795 => x"b387e700",
         796 => x"b3871741",
         797 => x"b3d8b702",
         798 => x"13180801",
         799 => x"13580801",
         800 => x"b3f7b702",
         801 => x"b3061603",
         802 => x"93970701",
         803 => x"3368f800",
         804 => x"93870800",
         805 => x"637cd800",
         806 => x"33080701",
         807 => x"9387f8ff",
         808 => x"6366e800",
         809 => x"6374d800",
         810 => x"9387e8ff",
         811 => x"13150501",
         812 => x"3365f500",
         813 => x"93050000",
         814 => x"67800000",
         815 => x"37050001",
         816 => x"93060001",
         817 => x"e36ca6f2",
         818 => x"93068001",
         819 => x"6ff01ff3",
         820 => x"63140600",
         821 => x"73001000",
         822 => x"b7070100",
         823 => x"6370f60c",
         824 => x"93360610",
         825 => x"93c61600",
         826 => x"93963600",
         827 => x"b357d600",
         828 => x"b385f500",
         829 => x"83c70500",
         830 => x"b387d700",
         831 => x"93060002",
         832 => x"b385f640",
         833 => x"6396f60a",
         834 => x"b387c840",
         835 => x"93051000",
         836 => x"93580701",
         837 => x"33de1703",
         838 => x"13160701",
         839 => x"13560601",
         840 => x"93560801",
         841 => x"b3f71703",
         842 => x"13050e00",
         843 => x"3303c603",
         844 => x"93970701",
         845 => x"b3e7f600",
         846 => x"63fe6700",
         847 => x"b387e700",
         848 => x"1305feff",
         849 => x"63e8e700",
         850 => x"63f66700",
         851 => x"1305eeff",
         852 => x"b387e700",
         853 => x"b3876740",
         854 => x"33d31703",
         855 => x"13180801",
         856 => x"13580801",
         857 => x"b3f71703",
         858 => x"b3066602",
         859 => x"93970701",
         860 => x"3368f800",
         861 => x"93070300",
         862 => x"637cd800",
         863 => x"33080701",
         864 => x"9307f3ff",
         865 => x"6366e800",
         866 => x"6374d800",
         867 => x"9307e3ff",
         868 => x"13150501",
         869 => x"3365f500",
         870 => x"67800000",
         871 => x"b7070001",
         872 => x"93060001",
         873 => x"e364f6f4",
         874 => x"93068001",
         875 => x"6ff01ff4",
         876 => x"3317b600",
         877 => x"b3d6f800",
         878 => x"13550701",
         879 => x"b357f300",
         880 => x"3318b300",
         881 => x"33d3a602",
         882 => x"13160701",
         883 => x"b398b800",
         884 => x"13560601",
         885 => x"b3e71701",
         886 => x"b3f6a602",
         887 => x"b3086602",
         888 => x"93950601",
         889 => x"93d60701",
         890 => x"b3e6b600",
         891 => x"93050300",
         892 => x"63fe1601",
         893 => x"b386e600",
         894 => x"9305f3ff",
         895 => x"63e8e600",
         896 => x"63f61601",
         897 => x"9305e3ff",
         898 => x"b386e600",
         899 => x"b3861641",
         900 => x"b3d8a602",
         901 => x"93970701",
         902 => x"93d70701",
         903 => x"b3f6a602",
         904 => x"33061603",
         905 => x"93960601",
         906 => x"b3e7d700",
         907 => x"93860800",
         908 => x"63fec700",
         909 => x"b387e700",
         910 => x"9386f8ff",
         911 => x"63e8e700",
         912 => x"63f6c700",
         913 => x"9386e8ff",
         914 => x"b387e700",
         915 => x"93950501",
         916 => x"b387c740",
         917 => x"b3e5d500",
         918 => x"6ff09feb",
         919 => x"63e6d518",
         920 => x"b7070100",
         921 => x"63f4f604",
         922 => x"13b70610",
         923 => x"13471700",
         924 => x"13173700",
         925 => x"b7370000",
         926 => x"b3d5e600",
         927 => x"9387c7d2",
         928 => x"b387b700",
         929 => x"83c70700",
         930 => x"b387e700",
         931 => x"13070002",
         932 => x"b305f740",
         933 => x"6316f702",
         934 => x"13051000",
         935 => x"e3ee16e1",
         936 => x"3335c300",
         937 => x"13451500",
         938 => x"67800000",
         939 => x"b7070001",
         940 => x"13070001",
         941 => x"e3e0f6fc",
         942 => x"13078001",
         943 => x"6ff09ffb",
         944 => x"3357f600",
         945 => x"b396b600",
         946 => x"b366d700",
         947 => x"33d7f800",
         948 => x"b398b800",
         949 => x"b357f300",
         950 => x"b3e71701",
         951 => x"93d80601",
         952 => x"b35e1703",
         953 => x"13980601",
         954 => x"13580801",
         955 => x"3316b600",
         956 => x"33771703",
         957 => x"330ed803",
         958 => x"13150701",
         959 => x"13d70701",
         960 => x"3367a700",
         961 => x"13850e00",
         962 => x"637ec701",
         963 => x"3307d700",
         964 => x"1385feff",
         965 => x"6368d700",
         966 => x"6376c701",
         967 => x"1385eeff",
         968 => x"3307d700",
         969 => x"3307c741",
         970 => x"335e1703",
         971 => x"93970701",
         972 => x"93d70701",
         973 => x"33771703",
         974 => x"3308c803",
         975 => x"13170701",
         976 => x"b3e7e700",
         977 => x"13070e00",
         978 => x"63fe0701",
         979 => x"b387d700",
         980 => x"1307feff",
         981 => x"63e8d700",
         982 => x"63f60701",
         983 => x"1307eeff",
         984 => x"b387d700",
         985 => x"13150501",
         986 => x"370e0100",
         987 => x"3365e500",
         988 => x"9306feff",
         989 => x"3377d500",
         990 => x"b3870741",
         991 => x"b376d600",
         992 => x"13580501",
         993 => x"13560601",
         994 => x"b308d702",
         995 => x"b306d802",
         996 => x"3307c702",
         997 => x"3308c802",
         998 => x"3306d700",
         999 => x"13d70801",
        1000 => x"3307c700",
        1001 => x"6374d700",
        1002 => x"3308c801",
        1003 => x"93560701",
        1004 => x"b3860601",
        1005 => x"63e6d702",
        1006 => x"e39ed7ce",
        1007 => x"b7070100",
        1008 => x"9387f7ff",
        1009 => x"3377f700",
        1010 => x"13170701",
        1011 => x"b3f8f800",
        1012 => x"3313b300",
        1013 => x"33071701",
        1014 => x"93050000",
        1015 => x"e37ee3cc",
        1016 => x"1305f5ff",
        1017 => x"6ff01fcd",
        1018 => x"93050000",
        1019 => x"13050000",
        1020 => x"67800000",
        1021 => x"13080600",
        1022 => x"93070500",
        1023 => x"13870500",
        1024 => x"63960620",
        1025 => x"b7380000",
        1026 => x"9388c8d2",
        1027 => x"63fcc50c",
        1028 => x"b7060100",
        1029 => x"637ed60a",
        1030 => x"93360610",
        1031 => x"93c61600",
        1032 => x"93963600",
        1033 => x"3353d600",
        1034 => x"b3886800",
        1035 => x"83c80800",
        1036 => x"13030002",
        1037 => x"b386d800",
        1038 => x"b308d340",
        1039 => x"630cd300",
        1040 => x"33971501",
        1041 => x"b356d500",
        1042 => x"33181601",
        1043 => x"33e7e600",
        1044 => x"b3171501",
        1045 => x"13560801",
        1046 => x"b356c702",
        1047 => x"13150801",
        1048 => x"13550501",
        1049 => x"3377c702",
        1050 => x"b386a602",
        1051 => x"93150701",
        1052 => x"13d70701",
        1053 => x"3367b700",
        1054 => x"637ad700",
        1055 => x"33070701",
        1056 => x"63660701",
        1057 => x"6374d700",
        1058 => x"33070701",
        1059 => x"3307d740",
        1060 => x"b356c702",
        1061 => x"3377c702",
        1062 => x"b386a602",
        1063 => x"93970701",
        1064 => x"13170701",
        1065 => x"93d70701",
        1066 => x"b3e7e700",
        1067 => x"63fad700",
        1068 => x"b3870701",
        1069 => x"63e60701",
        1070 => x"63f4d700",
        1071 => x"b3870701",
        1072 => x"b387d740",
        1073 => x"33d51701",
        1074 => x"93050000",
        1075 => x"67800000",
        1076 => x"37030001",
        1077 => x"93060001",
        1078 => x"e36666f4",
        1079 => x"93068001",
        1080 => x"6ff05ff4",
        1081 => x"63140600",
        1082 => x"73001000",
        1083 => x"37070100",
        1084 => x"637ee606",
        1085 => x"93360610",
        1086 => x"93c61600",
        1087 => x"93963600",
        1088 => x"3357d600",
        1089 => x"b388e800",
        1090 => x"03c70800",
        1091 => x"3307d700",
        1092 => x"93060002",
        1093 => x"b388e640",
        1094 => x"6394e606",
        1095 => x"3387c540",
        1096 => x"93550801",
        1097 => x"3356b702",
        1098 => x"13150801",
        1099 => x"13550501",
        1100 => x"93d60701",
        1101 => x"3377b702",
        1102 => x"3306a602",
        1103 => x"13170701",
        1104 => x"33e7e600",
        1105 => x"637ac700",
        1106 => x"33070701",
        1107 => x"63660701",
        1108 => x"6374c700",
        1109 => x"33070701",
        1110 => x"3307c740",
        1111 => x"b356b702",
        1112 => x"3377b702",
        1113 => x"b386a602",
        1114 => x"6ff05ff3",
        1115 => x"37070001",
        1116 => x"93060001",
        1117 => x"e366e6f8",
        1118 => x"93068001",
        1119 => x"6ff05ff8",
        1120 => x"33181601",
        1121 => x"b3d6e500",
        1122 => x"b3171501",
        1123 => x"b3951501",
        1124 => x"3357e500",
        1125 => x"13550801",
        1126 => x"3367b700",
        1127 => x"b3d5a602",
        1128 => x"13130801",
        1129 => x"13530301",
        1130 => x"b3f6a602",
        1131 => x"b3856502",
        1132 => x"13960601",
        1133 => x"93560701",
        1134 => x"b3e6c600",
        1135 => x"63fab600",
        1136 => x"b3860601",
        1137 => x"63e60601",
        1138 => x"63f4b600",
        1139 => x"b3860601",
        1140 => x"b386b640",
        1141 => x"33d6a602",
        1142 => x"13170701",
        1143 => x"13570701",
        1144 => x"b3f6a602",
        1145 => x"33066602",
        1146 => x"93960601",
        1147 => x"3367d700",
        1148 => x"637ac700",
        1149 => x"33070701",
        1150 => x"63660701",
        1151 => x"6374c700",
        1152 => x"33070701",
        1153 => x"3307c740",
        1154 => x"6ff09ff1",
        1155 => x"63e4d51c",
        1156 => x"37080100",
        1157 => x"63fe0605",
        1158 => x"13b80610",
        1159 => x"13481800",
        1160 => x"13183800",
        1161 => x"b7380000",
        1162 => x"33d30601",
        1163 => x"9388c8d2",
        1164 => x"b3886800",
        1165 => x"83c80800",
        1166 => x"13030002",
        1167 => x"b3880801",
        1168 => x"33081341",
        1169 => x"63101305",
        1170 => x"63e4b600",
        1171 => x"636cc500",
        1172 => x"3306c540",
        1173 => x"b386d540",
        1174 => x"3337c500",
        1175 => x"3387e640",
        1176 => x"93070600",
        1177 => x"13850700",
        1178 => x"93050700",
        1179 => x"67800000",
        1180 => x"b7080001",
        1181 => x"13080001",
        1182 => x"e3e616fb",
        1183 => x"13088001",
        1184 => x"6ff05ffa",
        1185 => x"b3960601",
        1186 => x"33531601",
        1187 => x"3363d300",
        1188 => x"135e0301",
        1189 => x"b3d61501",
        1190 => x"33dfc603",
        1191 => x"13170301",
        1192 => x"13570701",
        1193 => x"b3970501",
        1194 => x"b3551501",
        1195 => x"b3e5f500",
        1196 => x"93d70501",
        1197 => x"33160601",
        1198 => x"33150501",
        1199 => x"b3f6c603",
        1200 => x"b30ee703",
        1201 => x"93960601",
        1202 => x"b3e7d700",
        1203 => x"93060f00",
        1204 => x"63fed701",
        1205 => x"b3876700",
        1206 => x"9306ffff",
        1207 => x"63e86700",
        1208 => x"63f6d701",
        1209 => x"9306efff",
        1210 => x"b3876700",
        1211 => x"b387d741",
        1212 => x"b3dec703",
        1213 => x"93950501",
        1214 => x"93d50501",
        1215 => x"b3f7c703",
        1216 => x"3307d703",
        1217 => x"93970701",
        1218 => x"b3e5f500",
        1219 => x"93870e00",
        1220 => x"63fee500",
        1221 => x"b3856500",
        1222 => x"9387feff",
        1223 => x"63e86500",
        1224 => x"63f6e500",
        1225 => x"9387eeff",
        1226 => x"b3856500",
        1227 => x"93960601",
        1228 => x"370f0100",
        1229 => x"b3e6f600",
        1230 => x"9307ffff",
        1231 => x"135e0601",
        1232 => x"b385e540",
        1233 => x"33f7f600",
        1234 => x"93d60601",
        1235 => x"b377f600",
        1236 => x"b30ef702",
        1237 => x"b387f602",
        1238 => x"3307c703",
        1239 => x"b386c603",
        1240 => x"330ef700",
        1241 => x"13d70e01",
        1242 => x"3307c701",
        1243 => x"6374f700",
        1244 => x"b386e601",
        1245 => x"93570701",
        1246 => x"b387d700",
        1247 => x"b7060100",
        1248 => x"9386f6ff",
        1249 => x"3377d700",
        1250 => x"13170701",
        1251 => x"b3fede00",
        1252 => x"3307d701",
        1253 => x"63e6f500",
        1254 => x"639ef500",
        1255 => x"637ce500",
        1256 => x"3306c740",
        1257 => x"3337c700",
        1258 => x"33076700",
        1259 => x"b387e740",
        1260 => x"13070600",
        1261 => x"3307e540",
        1262 => x"3335e500",
        1263 => x"b385f540",
        1264 => x"b385a540",
        1265 => x"b3981501",
        1266 => x"33570701",
        1267 => x"33e5e800",
        1268 => x"b3d50501",
        1269 => x"67800000",
        1270 => x"13030500",
        1271 => x"630e0600",
        1272 => x"83830500",
        1273 => x"23007300",
        1274 => x"1306f6ff",
        1275 => x"13031300",
        1276 => x"93851500",
        1277 => x"e31606fe",
        1278 => x"67800000",
        1279 => x"13030500",
        1280 => x"630a0600",
        1281 => x"2300b300",
        1282 => x"1306f6ff",
        1283 => x"13031300",
        1284 => x"e31a06fe",
        1285 => x"67800000",
        1286 => x"630c0602",
        1287 => x"13030500",
        1288 => x"93061000",
        1289 => x"636ab500",
        1290 => x"9306f0ff",
        1291 => x"1307f6ff",
        1292 => x"3303e300",
        1293 => x"b385e500",
        1294 => x"83830500",
        1295 => x"23007300",
        1296 => x"1306f6ff",
        1297 => x"3303d300",
        1298 => x"b385d500",
        1299 => x"e31606fe",
        1300 => x"67800000",
        1301 => x"130101f8",
        1302 => x"232c8106",
        1303 => x"23263107",
        1304 => x"232e1106",
        1305 => x"232a9106",
        1306 => x"23282107",
        1307 => x"23244107",
        1308 => x"23225107",
        1309 => x"23206107",
        1310 => x"232e7105",
        1311 => x"232c8105",
        1312 => x"232a9105",
        1313 => x"2328a105",
        1314 => x"2326b105",
        1315 => x"93090500",
        1316 => x"13840500",
        1317 => x"232c0100",
        1318 => x"232e0100",
        1319 => x"23200102",
        1320 => x"23220102",
        1321 => x"23240102",
        1322 => x"23260102",
        1323 => x"23280102",
        1324 => x"232a0102",
        1325 => x"232c0102",
        1326 => x"232e0102",
        1327 => x"97f2ffff",
        1328 => x"938282e1",
        1329 => x"73905230",
        1330 => x"efe05fbb",
        1331 => x"b7877d01",
        1332 => x"370700f0",
        1333 => x"9387f783",
        1334 => x"2326f708",
        1335 => x"93071001",
        1336 => x"2320f708",
        1337 => x"b7220000",
        1338 => x"93828280",
        1339 => x"73900230",
        1340 => x"37390000",
        1341 => x"130589e5",
        1342 => x"efe01fbc",
        1343 => x"63543003",
        1344 => x"9384f9ff",
        1345 => x"9309f0ff",
        1346 => x"03250400",
        1347 => x"9384f4ff",
        1348 => x"13044400",
        1349 => x"efe05fba",
        1350 => x"130589e5",
        1351 => x"efe0dfb9",
        1352 => x"e39434ff",
        1353 => x"37350000",
        1354 => x"b7faeeee",
        1355 => x"1305c5e2",
        1356 => x"b7040010",
        1357 => x"37190000",
        1358 => x"1384faee",
        1359 => x"efe0dfb7",
        1360 => x"130c0000",
        1361 => x"b73b0000",
        1362 => x"9384f4ff",
        1363 => x"130bf000",
        1364 => x"938aeaee",
        1365 => x"130909e1",
        1366 => x"93090000",
        1367 => x"130a0019",
        1368 => x"93050000",
        1369 => x"13058100",
        1370 => x"ef008035",
        1371 => x"130c1c00",
        1372 => x"63020502",
        1373 => x"e3164cff",
        1374 => x"73001000",
        1375 => x"93050000",
        1376 => x"13058100",
        1377 => x"130c0000",
        1378 => x"ef008033",
        1379 => x"130c1c00",
        1380 => x"e31205fe",
        1381 => x"832c8100",
        1382 => x"8325c100",
        1383 => x"13060900",
        1384 => x"93d7cc01",
        1385 => x"13974500",
        1386 => x"b367f700",
        1387 => x"b3f79700",
        1388 => x"33f79c00",
        1389 => x"13d5f541",
        1390 => x"13d88501",
        1391 => x"3307f700",
        1392 => x"33070701",
        1393 => x"9377d500",
        1394 => x"3307f700",
        1395 => x"33776703",
        1396 => x"937725ff",
        1397 => x"93860900",
        1398 => x"13850c00",
        1399 => x"3307f700",
        1400 => x"b387ec40",
        1401 => x"1357f741",
        1402 => x"33b8fc00",
        1403 => x"3387e540",
        1404 => x"33070741",
        1405 => x"b3885703",
        1406 => x"33078702",
        1407 => x"33b88702",
        1408 => x"33071701",
        1409 => x"b3878702",
        1410 => x"33070701",
        1411 => x"1358f741",
        1412 => x"13783800",
        1413 => x"b307f800",
        1414 => x"33b80701",
        1415 => x"3307e800",
        1416 => x"1318e701",
        1417 => x"93d72700",
        1418 => x"b367f800",
        1419 => x"93582740",
        1420 => x"13984800",
        1421 => x"13d3c701",
        1422 => x"33636800",
        1423 => x"33739300",
        1424 => x"33f89700",
        1425 => x"13de8801",
        1426 => x"1357f741",
        1427 => x"33086800",
        1428 => x"3308c801",
        1429 => x"1373d700",
        1430 => x"33086800",
        1431 => x"33786803",
        1432 => x"137727ff",
        1433 => x"139d4700",
        1434 => x"330dfd40",
        1435 => x"131d2d00",
        1436 => x"338dac41",
        1437 => x"3308e800",
        1438 => x"33870741",
        1439 => x"1358f841",
        1440 => x"33b3e700",
        1441 => x"b3880841",
        1442 => x"b3886840",
        1443 => x"b3888802",
        1444 => x"33035703",
        1445 => x"33388702",
        1446 => x"b3886800",
        1447 => x"33078702",
        1448 => x"b3880801",
        1449 => x"13d8f841",
        1450 => x"13783800",
        1451 => x"3307e800",
        1452 => x"33380701",
        1453 => x"33081801",
        1454 => x"1318e801",
        1455 => x"13572700",
        1456 => x"3367e800",
        1457 => x"13184700",
        1458 => x"3307e840",
        1459 => x"13172700",
        1460 => x"b38de740",
        1461 => x"eff08f87",
        1462 => x"83260101",
        1463 => x"13070500",
        1464 => x"13080d00",
        1465 => x"93870d00",
        1466 => x"13860c00",
        1467 => x"9385cbe5",
        1468 => x"13058101",
        1469 => x"ef00c015",
        1470 => x"13058101",
        1471 => x"efe0df9b",
        1472 => x"e3104ce7",
        1473 => x"6ff05fe7",
        1474 => x"03a5c187",
        1475 => x"67800000",
        1476 => x"130101ff",
        1477 => x"23248100",
        1478 => x"23261100",
        1479 => x"93070000",
        1480 => x"13040500",
        1481 => x"63880700",
        1482 => x"93050000",
        1483 => x"97000000",
        1484 => x"e7000000",
        1485 => x"b7370000",
        1486 => x"03a547fd",
        1487 => x"83278502",
        1488 => x"63840700",
        1489 => x"e7800700",
        1490 => x"13050400",
        1491 => x"ef108033",
        1492 => x"130101ff",
        1493 => x"23248100",
        1494 => x"23229100",
        1495 => x"37340000",
        1496 => x"b7340000",
        1497 => x"938784fd",
        1498 => x"130484fd",
        1499 => x"3304f440",
        1500 => x"23202101",
        1501 => x"23261100",
        1502 => x"13542440",
        1503 => x"938484fd",
        1504 => x"13090000",
        1505 => x"63108904",
        1506 => x"b7340000",
        1507 => x"37340000",
        1508 => x"938784fd",
        1509 => x"130484fd",
        1510 => x"3304f440",
        1511 => x"13542440",
        1512 => x"938484fd",
        1513 => x"13090000",
        1514 => x"63188902",
        1515 => x"8320c100",
        1516 => x"03248100",
        1517 => x"83244100",
        1518 => x"03290100",
        1519 => x"13010101",
        1520 => x"67800000",
        1521 => x"83a70400",
        1522 => x"13091900",
        1523 => x"93844400",
        1524 => x"e7800700",
        1525 => x"6ff01ffb",
        1526 => x"83a70400",
        1527 => x"13091900",
        1528 => x"93844400",
        1529 => x"e7800700",
        1530 => x"6ff01ffc",
        1531 => x"130101f6",
        1532 => x"232af108",
        1533 => x"b7070080",
        1534 => x"93c7f7ff",
        1535 => x"232ef100",
        1536 => x"2328f100",
        1537 => x"b707ffff",
        1538 => x"2326d108",
        1539 => x"2324b100",
        1540 => x"232cb100",
        1541 => x"93878720",
        1542 => x"9306c108",
        1543 => x"93058100",
        1544 => x"232e1106",
        1545 => x"232af100",
        1546 => x"2328e108",
        1547 => x"232c0109",
        1548 => x"232e1109",
        1549 => x"2322d100",
        1550 => x"ef004041",
        1551 => x"83278100",
        1552 => x"23800700",
        1553 => x"8320c107",
        1554 => x"1301010a",
        1555 => x"67800000",
        1556 => x"130101f6",
        1557 => x"232af108",
        1558 => x"b7070080",
        1559 => x"93c7f7ff",
        1560 => x"232ef100",
        1561 => x"2328f100",
        1562 => x"b707ffff",
        1563 => x"93878720",
        1564 => x"232af100",
        1565 => x"2324a100",
        1566 => x"232ca100",
        1567 => x"03a5c187",
        1568 => x"2324c108",
        1569 => x"2326d108",
        1570 => x"13860500",
        1571 => x"93068108",
        1572 => x"93058100",
        1573 => x"232e1106",
        1574 => x"2328e108",
        1575 => x"232c0109",
        1576 => x"232e1109",
        1577 => x"2322d100",
        1578 => x"ef00403a",
        1579 => x"83278100",
        1580 => x"23800700",
        1581 => x"8320c107",
        1582 => x"1301010a",
        1583 => x"67800000",
        1584 => x"13860500",
        1585 => x"93050500",
        1586 => x"03a5c187",
        1587 => x"6f004000",
        1588 => x"130101ff",
        1589 => x"23248100",
        1590 => x"23229100",
        1591 => x"13040500",
        1592 => x"13850500",
        1593 => x"93050600",
        1594 => x"23261100",
        1595 => x"23a20188",
        1596 => x"ef10401c",
        1597 => x"9307f0ff",
        1598 => x"6318f500",
        1599 => x"83a74188",
        1600 => x"63840700",
        1601 => x"2320f400",
        1602 => x"8320c100",
        1603 => x"03248100",
        1604 => x"83244100",
        1605 => x"13010101",
        1606 => x"67800000",
        1607 => x"130101fe",
        1608 => x"23282101",
        1609 => x"03a98500",
        1610 => x"232c8100",
        1611 => x"23263101",
        1612 => x"23244101",
        1613 => x"23225101",
        1614 => x"232e1100",
        1615 => x"232a9100",
        1616 => x"23206101",
        1617 => x"83aa0500",
        1618 => x"13840500",
        1619 => x"130a0600",
        1620 => x"93890600",
        1621 => x"63ec2609",
        1622 => x"83d7c500",
        1623 => x"13f70748",
        1624 => x"63040708",
        1625 => x"03274401",
        1626 => x"93043000",
        1627 => x"83a50501",
        1628 => x"b384e402",
        1629 => x"13072000",
        1630 => x"b38aba40",
        1631 => x"130b0500",
        1632 => x"b3c4e402",
        1633 => x"13871600",
        1634 => x"33075701",
        1635 => x"63f4e400",
        1636 => x"93040700",
        1637 => x"93f70740",
        1638 => x"6386070a",
        1639 => x"93850400",
        1640 => x"13050b00",
        1641 => x"ef001065",
        1642 => x"13090500",
        1643 => x"630c050a",
        1644 => x"83250401",
        1645 => x"13860a00",
        1646 => x"eff01fa2",
        1647 => x"8357c400",
        1648 => x"93f7f7b7",
        1649 => x"93e70708",
        1650 => x"2316f400",
        1651 => x"23282401",
        1652 => x"232a9400",
        1653 => x"33095901",
        1654 => x"b3845441",
        1655 => x"23202401",
        1656 => x"23249400",
        1657 => x"13890900",
        1658 => x"63f42901",
        1659 => x"13890900",
        1660 => x"03250400",
        1661 => x"13060900",
        1662 => x"93050a00",
        1663 => x"eff0dfa1",
        1664 => x"83278400",
        1665 => x"13050000",
        1666 => x"b3872741",
        1667 => x"2324f400",
        1668 => x"83270400",
        1669 => x"b3872701",
        1670 => x"2320f400",
        1671 => x"8320c101",
        1672 => x"03248101",
        1673 => x"83244101",
        1674 => x"03290101",
        1675 => x"8329c100",
        1676 => x"032a8100",
        1677 => x"832a4100",
        1678 => x"032b0100",
        1679 => x"13010102",
        1680 => x"67800000",
        1681 => x"13860400",
        1682 => x"13050b00",
        1683 => x"ef00906f",
        1684 => x"13090500",
        1685 => x"e31c05f6",
        1686 => x"83250401",
        1687 => x"13050b00",
        1688 => x"ef00d049",
        1689 => x"9307c000",
        1690 => x"2320fb00",
        1691 => x"8357c400",
        1692 => x"1305f0ff",
        1693 => x"93e70704",
        1694 => x"2316f400",
        1695 => x"6ff01ffa",
        1696 => x"83278600",
        1697 => x"130101fd",
        1698 => x"232e3101",
        1699 => x"23286101",
        1700 => x"23261102",
        1701 => x"23248102",
        1702 => x"23229102",
        1703 => x"23202103",
        1704 => x"232c4101",
        1705 => x"232a5101",
        1706 => x"23267101",
        1707 => x"23248101",
        1708 => x"23229101",
        1709 => x"2320a101",
        1710 => x"032b0600",
        1711 => x"93090600",
        1712 => x"63980712",
        1713 => x"13050000",
        1714 => x"8320c102",
        1715 => x"03248102",
        1716 => x"23a20900",
        1717 => x"83244102",
        1718 => x"03290102",
        1719 => x"8329c101",
        1720 => x"032a8101",
        1721 => x"832a4101",
        1722 => x"032b0101",
        1723 => x"832bc100",
        1724 => x"032c8100",
        1725 => x"832c4100",
        1726 => x"032d0100",
        1727 => x"13010103",
        1728 => x"67800000",
        1729 => x"832a0b00",
        1730 => x"032d4b00",
        1731 => x"130b8b00",
        1732 => x"03298400",
        1733 => x"832c0400",
        1734 => x"e3060dfe",
        1735 => x"63642d09",
        1736 => x"8357c400",
        1737 => x"13f70748",
        1738 => x"630e0706",
        1739 => x"83244401",
        1740 => x"83250401",
        1741 => x"b3849b02",
        1742 => x"b38cbc40",
        1743 => x"13871c00",
        1744 => x"3307a701",
        1745 => x"b3c48403",
        1746 => x"63f4e400",
        1747 => x"93040700",
        1748 => x"93f70740",
        1749 => x"638c070a",
        1750 => x"93850400",
        1751 => x"13050a00",
        1752 => x"ef005049",
        1753 => x"13090500",
        1754 => x"6302050c",
        1755 => x"83250401",
        1756 => x"13860c00",
        1757 => x"eff05f86",
        1758 => x"8357c400",
        1759 => x"93f7f7b7",
        1760 => x"93e70708",
        1761 => x"2316f400",
        1762 => x"23282401",
        1763 => x"232a9400",
        1764 => x"33099901",
        1765 => x"b3849441",
        1766 => x"23202401",
        1767 => x"23249400",
        1768 => x"13090d00",
        1769 => x"63742d01",
        1770 => x"13090d00",
        1771 => x"03250400",
        1772 => x"93850a00",
        1773 => x"13060900",
        1774 => x"eff01f86",
        1775 => x"83278400",
        1776 => x"b38aaa01",
        1777 => x"b3872741",
        1778 => x"2324f400",
        1779 => x"83270400",
        1780 => x"b3872701",
        1781 => x"2320f400",
        1782 => x"83a78900",
        1783 => x"b387a741",
        1784 => x"23a4f900",
        1785 => x"e38007ee",
        1786 => x"130d0000",
        1787 => x"6ff05ff2",
        1788 => x"130a0500",
        1789 => x"13840500",
        1790 => x"930a0000",
        1791 => x"130d0000",
        1792 => x"930b3000",
        1793 => x"130c2000",
        1794 => x"6ff09ff0",
        1795 => x"13860400",
        1796 => x"13050a00",
        1797 => x"ef001053",
        1798 => x"13090500",
        1799 => x"e31605f6",
        1800 => x"83250401",
        1801 => x"13050a00",
        1802 => x"ef00502d",
        1803 => x"9307c000",
        1804 => x"2320fa00",
        1805 => x"8357c400",
        1806 => x"1305f0ff",
        1807 => x"93e70704",
        1808 => x"2316f400",
        1809 => x"23a40900",
        1810 => x"6ff01fe8",
        1811 => x"83d7c500",
        1812 => x"130101f5",
        1813 => x"2324810a",
        1814 => x"2322910a",
        1815 => x"2320210b",
        1816 => x"232c4109",
        1817 => x"2326110a",
        1818 => x"232e3109",
        1819 => x"232a5109",
        1820 => x"23286109",
        1821 => x"23267109",
        1822 => x"23248109",
        1823 => x"23229109",
        1824 => x"2320a109",
        1825 => x"232eb107",
        1826 => x"93f70708",
        1827 => x"130a0500",
        1828 => x"13890500",
        1829 => x"93040600",
        1830 => x"13840600",
        1831 => x"63880706",
        1832 => x"83a70501",
        1833 => x"63940706",
        1834 => x"93050004",
        1835 => x"ef009034",
        1836 => x"2320a900",
        1837 => x"2328a900",
        1838 => x"63160504",
        1839 => x"9307c000",
        1840 => x"2320fa00",
        1841 => x"1305f0ff",
        1842 => x"8320c10a",
        1843 => x"0324810a",
        1844 => x"8324410a",
        1845 => x"0329010a",
        1846 => x"8329c109",
        1847 => x"032a8109",
        1848 => x"832a4109",
        1849 => x"032b0109",
        1850 => x"832bc108",
        1851 => x"032c8108",
        1852 => x"832c4108",
        1853 => x"032d0108",
        1854 => x"832dc107",
        1855 => x"1301010b",
        1856 => x"67800000",
        1857 => x"93070004",
        1858 => x"232af900",
        1859 => x"93070002",
        1860 => x"a304f102",
        1861 => x"93070003",
        1862 => x"23220102",
        1863 => x"2305f102",
        1864 => x"23268100",
        1865 => x"930c5002",
        1866 => x"373b0000",
        1867 => x"b73b0000",
        1868 => x"373d0000",
        1869 => x"372c0000",
        1870 => x"930a0000",
        1871 => x"13840400",
        1872 => x"83470400",
        1873 => x"63840700",
        1874 => x"639c970d",
        1875 => x"b30d9440",
        1876 => x"63069402",
        1877 => x"93860d00",
        1878 => x"13860400",
        1879 => x"93050900",
        1880 => x"13050a00",
        1881 => x"eff09fbb",
        1882 => x"9307f0ff",
        1883 => x"6306f524",
        1884 => x"83274102",
        1885 => x"b387b701",
        1886 => x"2322f102",
        1887 => x"83470400",
        1888 => x"638c0722",
        1889 => x"9307f0ff",
        1890 => x"93041400",
        1891 => x"23280100",
        1892 => x"232e0100",
        1893 => x"232af100",
        1894 => x"232c0100",
        1895 => x"a3090104",
        1896 => x"23240106",
        1897 => x"930d1000",
        1898 => x"83c50400",
        1899 => x"13065000",
        1900 => x"13050bf4",
        1901 => x"ef005012",
        1902 => x"83270101",
        1903 => x"13841400",
        1904 => x"63140506",
        1905 => x"13f70701",
        1906 => x"63060700",
        1907 => x"13070002",
        1908 => x"a309e104",
        1909 => x"13f78700",
        1910 => x"63060700",
        1911 => x"1307b002",
        1912 => x"a309e104",
        1913 => x"83c60400",
        1914 => x"1307a002",
        1915 => x"638ce604",
        1916 => x"8327c101",
        1917 => x"13840400",
        1918 => x"93060000",
        1919 => x"13069000",
        1920 => x"1305a000",
        1921 => x"03470400",
        1922 => x"93051400",
        1923 => x"130707fd",
        1924 => x"637ce608",
        1925 => x"63840604",
        1926 => x"232ef100",
        1927 => x"6f000004",
        1928 => x"13041400",
        1929 => x"6ff0dff1",
        1930 => x"13070bf4",
        1931 => x"3305e540",
        1932 => x"3395ad00",
        1933 => x"b3e7a700",
        1934 => x"2328f100",
        1935 => x"93040400",
        1936 => x"6ff09ff6",
        1937 => x"0327c100",
        1938 => x"93064700",
        1939 => x"03270700",
        1940 => x"2326d100",
        1941 => x"63400704",
        1942 => x"232ee100",
        1943 => x"03470400",
        1944 => x"9307e002",
        1945 => x"6316f708",
        1946 => x"03471400",
        1947 => x"9307a002",
        1948 => x"631af704",
        1949 => x"8327c100",
        1950 => x"13042400",
        1951 => x"13874700",
        1952 => x"83a70700",
        1953 => x"2326e100",
        1954 => x"63ca0702",
        1955 => x"232af100",
        1956 => x"6f000006",
        1957 => x"3307e040",
        1958 => x"93e72700",
        1959 => x"232ee100",
        1960 => x"2328f100",
        1961 => x"6ff09ffb",
        1962 => x"b387a702",
        1963 => x"13840500",
        1964 => x"93061000",
        1965 => x"b387e700",
        1966 => x"6ff0dff4",
        1967 => x"9307f0ff",
        1968 => x"6ff0dffc",
        1969 => x"13041400",
        1970 => x"232a0100",
        1971 => x"93060000",
        1972 => x"93070000",
        1973 => x"13069000",
        1974 => x"1305a000",
        1975 => x"03470400",
        1976 => x"93051400",
        1977 => x"130707fd",
        1978 => x"6372e608",
        1979 => x"e39006fa",
        1980 => x"83450400",
        1981 => x"13063000",
        1982 => x"13858bf4",
        1983 => x"ef00c07d",
        1984 => x"63020502",
        1985 => x"93878bf4",
        1986 => x"3305f540",
        1987 => x"83270101",
        1988 => x"13070004",
        1989 => x"3317a700",
        1990 => x"b3e7e700",
        1991 => x"13041400",
        1992 => x"2328f100",
        1993 => x"83450400",
        1994 => x"13066000",
        1995 => x"1305cdf4",
        1996 => x"93041400",
        1997 => x"2304b102",
        1998 => x"ef00007a",
        1999 => x"630a0508",
        2000 => x"63980a04",
        2001 => x"03270101",
        2002 => x"8327c100",
        2003 => x"13770710",
        2004 => x"63080702",
        2005 => x"93874700",
        2006 => x"2326f100",
        2007 => x"83274102",
        2008 => x"b3873701",
        2009 => x"2322f102",
        2010 => x"6ff05fdd",
        2011 => x"b387a702",
        2012 => x"13840500",
        2013 => x"93061000",
        2014 => x"b387e700",
        2015 => x"6ff01ff6",
        2016 => x"93877700",
        2017 => x"93f787ff",
        2018 => x"93878700",
        2019 => x"6ff0dffc",
        2020 => x"1307c100",
        2021 => x"9306cc91",
        2022 => x"13060900",
        2023 => x"93050101",
        2024 => x"13050a00",
        2025 => x"97000000",
        2026 => x"e7000000",
        2027 => x"9307f0ff",
        2028 => x"93090500",
        2029 => x"e314f5fa",
        2030 => x"8357c900",
        2031 => x"1305f0ff",
        2032 => x"93f70704",
        2033 => x"e39207d0",
        2034 => x"03254102",
        2035 => x"6ff0dfcf",
        2036 => x"1307c100",
        2037 => x"9306cc91",
        2038 => x"13060900",
        2039 => x"93050101",
        2040 => x"13050a00",
        2041 => x"ef00801b",
        2042 => x"6ff05ffc",
        2043 => x"130101fd",
        2044 => x"232c4101",
        2045 => x"83a70501",
        2046 => x"130a0700",
        2047 => x"03a78500",
        2048 => x"23248102",
        2049 => x"23202103",
        2050 => x"232e3101",
        2051 => x"232a5101",
        2052 => x"23261102",
        2053 => x"23229102",
        2054 => x"23286101",
        2055 => x"23267101",
        2056 => x"93090500",
        2057 => x"13840500",
        2058 => x"13090600",
        2059 => x"938a0600",
        2060 => x"63d4e700",
        2061 => x"93070700",
        2062 => x"2320f900",
        2063 => x"03473404",
        2064 => x"63060700",
        2065 => x"93871700",
        2066 => x"2320f900",
        2067 => x"83270400",
        2068 => x"93f70702",
        2069 => x"63880700",
        2070 => x"83270900",
        2071 => x"93872700",
        2072 => x"2320f900",
        2073 => x"83240400",
        2074 => x"93f46400",
        2075 => x"639e0400",
        2076 => x"130b9401",
        2077 => x"930bf0ff",
        2078 => x"8327c400",
        2079 => x"03270900",
        2080 => x"b387e740",
        2081 => x"63c2f408",
        2082 => x"83473404",
        2083 => x"b336f000",
        2084 => x"83270400",
        2085 => x"93f70702",
        2086 => x"6390070c",
        2087 => x"13063404",
        2088 => x"93850a00",
        2089 => x"13850900",
        2090 => x"e7000a00",
        2091 => x"9307f0ff",
        2092 => x"6308f506",
        2093 => x"83270400",
        2094 => x"13074000",
        2095 => x"93040000",
        2096 => x"93f76700",
        2097 => x"639ce700",
        2098 => x"8324c400",
        2099 => x"83270900",
        2100 => x"b384f440",
        2101 => x"63d40400",
        2102 => x"93040000",
        2103 => x"83278400",
        2104 => x"03270401",
        2105 => x"6356f700",
        2106 => x"b387e740",
        2107 => x"b384f400",
        2108 => x"13090000",
        2109 => x"1304a401",
        2110 => x"130bf0ff",
        2111 => x"63902409",
        2112 => x"13050000",
        2113 => x"6f000002",
        2114 => x"93061000",
        2115 => x"13060b00",
        2116 => x"93850a00",
        2117 => x"13850900",
        2118 => x"e7000a00",
        2119 => x"631a7503",
        2120 => x"1305f0ff",
        2121 => x"8320c102",
        2122 => x"03248102",
        2123 => x"83244102",
        2124 => x"03290102",
        2125 => x"8329c101",
        2126 => x"032a8101",
        2127 => x"832a4101",
        2128 => x"032b0101",
        2129 => x"832bc100",
        2130 => x"13010103",
        2131 => x"67800000",
        2132 => x"93841400",
        2133 => x"6ff05ff2",
        2134 => x"3307d400",
        2135 => x"13060003",
        2136 => x"a301c704",
        2137 => x"03475404",
        2138 => x"93871600",
        2139 => x"b307f400",
        2140 => x"93862600",
        2141 => x"a381e704",
        2142 => x"6ff05ff2",
        2143 => x"93061000",
        2144 => x"13060400",
        2145 => x"93850a00",
        2146 => x"13850900",
        2147 => x"e7000a00",
        2148 => x"e30865f9",
        2149 => x"13091900",
        2150 => x"6ff05ff6",
        2151 => x"130101fd",
        2152 => x"23248102",
        2153 => x"23229102",
        2154 => x"23202103",
        2155 => x"232e3101",
        2156 => x"23261102",
        2157 => x"232c4101",
        2158 => x"232a5101",
        2159 => x"23286101",
        2160 => x"83c88501",
        2161 => x"93078007",
        2162 => x"93040500",
        2163 => x"13840500",
        2164 => x"13090600",
        2165 => x"93890600",
        2166 => x"63ee1701",
        2167 => x"93072006",
        2168 => x"93863504",
        2169 => x"63ee1701",
        2170 => x"63840828",
        2171 => x"93078005",
        2172 => x"6388f822",
        2173 => x"930a2404",
        2174 => x"23011405",
        2175 => x"6f004004",
        2176 => x"9387d8f9",
        2177 => x"93f7f70f",
        2178 => x"13065001",
        2179 => x"e364f6fe",
        2180 => x"37360000",
        2181 => x"93972700",
        2182 => x"1306c6f7",
        2183 => x"b387c700",
        2184 => x"83a70700",
        2185 => x"67800700",
        2186 => x"83270700",
        2187 => x"938a2504",
        2188 => x"93864700",
        2189 => x"83a70700",
        2190 => x"2320d700",
        2191 => x"2381f504",
        2192 => x"93071000",
        2193 => x"6f008026",
        2194 => x"83a70500",
        2195 => x"03250700",
        2196 => x"13f60708",
        2197 => x"93054500",
        2198 => x"63060602",
        2199 => x"83270500",
        2200 => x"2320b700",
        2201 => x"37380000",
        2202 => x"63d80700",
        2203 => x"1307d002",
        2204 => x"b307f040",
        2205 => x"a301e404",
        2206 => x"130848f5",
        2207 => x"1307a000",
        2208 => x"6f008006",
        2209 => x"13f60704",
        2210 => x"83270500",
        2211 => x"2320b700",
        2212 => x"e30a06fc",
        2213 => x"93970701",
        2214 => x"93d70741",
        2215 => x"6ff09ffc",
        2216 => x"03a60500",
        2217 => x"83270700",
        2218 => x"13750608",
        2219 => x"93854700",
        2220 => x"63080500",
        2221 => x"2320b700",
        2222 => x"83a70700",
        2223 => x"6f004001",
        2224 => x"13760604",
        2225 => x"2320b700",
        2226 => x"e30806fe",
        2227 => x"83d70700",
        2228 => x"37380000",
        2229 => x"1307f006",
        2230 => x"130848f5",
        2231 => x"6388e814",
        2232 => x"1307a000",
        2233 => x"a3010404",
        2234 => x"03264400",
        2235 => x"2324c400",
        2236 => x"63480600",
        2237 => x"83250400",
        2238 => x"93f5b5ff",
        2239 => x"2320b400",
        2240 => x"63960700",
        2241 => x"938a0600",
        2242 => x"63040602",
        2243 => x"938a0600",
        2244 => x"33f6e702",
        2245 => x"938afaff",
        2246 => x"3306c800",
        2247 => x"03460600",
        2248 => x"2380ca00",
        2249 => x"13860700",
        2250 => x"b3d7e702",
        2251 => x"e372e6fe",
        2252 => x"93078000",
        2253 => x"6314f702",
        2254 => x"83270400",
        2255 => x"93f71700",
        2256 => x"638e0700",
        2257 => x"03274400",
        2258 => x"83270401",
        2259 => x"63c8e700",
        2260 => x"93070003",
        2261 => x"a38ffafe",
        2262 => x"938afaff",
        2263 => x"b3865641",
        2264 => x"2328d400",
        2265 => x"13870900",
        2266 => x"93060900",
        2267 => x"1306c100",
        2268 => x"93050400",
        2269 => x"13850400",
        2270 => x"eff05fc7",
        2271 => x"130af0ff",
        2272 => x"631c4513",
        2273 => x"1305f0ff",
        2274 => x"8320c102",
        2275 => x"03248102",
        2276 => x"83244102",
        2277 => x"03290102",
        2278 => x"8329c101",
        2279 => x"032a8101",
        2280 => x"832a4101",
        2281 => x"032b0101",
        2282 => x"13010103",
        2283 => x"67800000",
        2284 => x"83a70500",
        2285 => x"93e70702",
        2286 => x"23a0f500",
        2287 => x"37380000",
        2288 => x"93088007",
        2289 => x"130888f6",
        2290 => x"a3021405",
        2291 => x"03260400",
        2292 => x"83250700",
        2293 => x"13750608",
        2294 => x"83a70500",
        2295 => x"93854500",
        2296 => x"631a0500",
        2297 => x"13750604",
        2298 => x"63060500",
        2299 => x"93970701",
        2300 => x"93d70701",
        2301 => x"2320b700",
        2302 => x"13771600",
        2303 => x"63060700",
        2304 => x"13660602",
        2305 => x"2320c400",
        2306 => x"13070001",
        2307 => x"e39c07ec",
        2308 => x"03260400",
        2309 => x"1376f6fd",
        2310 => x"2320c400",
        2311 => x"6ff09fec",
        2312 => x"37380000",
        2313 => x"130848f5",
        2314 => x"6ff01ffa",
        2315 => x"13078000",
        2316 => x"6ff05feb",
        2317 => x"03a60500",
        2318 => x"83270700",
        2319 => x"83a54501",
        2320 => x"13780608",
        2321 => x"13854700",
        2322 => x"630a0800",
        2323 => x"2320a700",
        2324 => x"83a70700",
        2325 => x"23a0b700",
        2326 => x"6f008001",
        2327 => x"2320a700",
        2328 => x"13760604",
        2329 => x"83a70700",
        2330 => x"e30606fe",
        2331 => x"2390b700",
        2332 => x"23280400",
        2333 => x"938a0600",
        2334 => x"6ff0dfee",
        2335 => x"83270700",
        2336 => x"03a64500",
        2337 => x"93050000",
        2338 => x"93864700",
        2339 => x"2320d700",
        2340 => x"83aa0700",
        2341 => x"13850a00",
        2342 => x"ef000024",
        2343 => x"63060500",
        2344 => x"33055541",
        2345 => x"2322a400",
        2346 => x"83274400",
        2347 => x"2328f400",
        2348 => x"a3010404",
        2349 => x"6ff01feb",
        2350 => x"83260401",
        2351 => x"13860a00",
        2352 => x"93050900",
        2353 => x"13850400",
        2354 => x"e7800900",
        2355 => x"e30c45eb",
        2356 => x"83270400",
        2357 => x"93f72700",
        2358 => x"63940704",
        2359 => x"8327c100",
        2360 => x"0325c400",
        2361 => x"e352f5ea",
        2362 => x"13850700",
        2363 => x"6ff0dfe9",
        2364 => x"93061000",
        2365 => x"13860a00",
        2366 => x"93050900",
        2367 => x"13850400",
        2368 => x"e7800900",
        2369 => x"e30065e9",
        2370 => x"130a1a00",
        2371 => x"8327c400",
        2372 => x"0327c100",
        2373 => x"b387e740",
        2374 => x"e34cfafc",
        2375 => x"6ff01ffc",
        2376 => x"130a0000",
        2377 => x"930a9401",
        2378 => x"130bf0ff",
        2379 => x"6ff01ffe",
        2380 => x"130101ff",
        2381 => x"23248100",
        2382 => x"13840500",
        2383 => x"83a50500",
        2384 => x"23229100",
        2385 => x"23261100",
        2386 => x"93040500",
        2387 => x"63840500",
        2388 => x"eff01ffe",
        2389 => x"93050400",
        2390 => x"03248100",
        2391 => x"8320c100",
        2392 => x"13850400",
        2393 => x"83244100",
        2394 => x"13010101",
        2395 => x"6f000019",
        2396 => x"83a7c187",
        2397 => x"6380a716",
        2398 => x"83274502",
        2399 => x"130101fe",
        2400 => x"232c8100",
        2401 => x"232e1100",
        2402 => x"232a9100",
        2403 => x"23282101",
        2404 => x"23263101",
        2405 => x"13040500",
        2406 => x"63840702",
        2407 => x"83a7c700",
        2408 => x"93040000",
        2409 => x"13090008",
        2410 => x"6392070e",
        2411 => x"83274402",
        2412 => x"83a50700",
        2413 => x"63860500",
        2414 => x"13050400",
        2415 => x"ef000014",
        2416 => x"83254401",
        2417 => x"63860500",
        2418 => x"13050400",
        2419 => x"ef000013",
        2420 => x"83254402",
        2421 => x"63860500",
        2422 => x"13050400",
        2423 => x"ef000012",
        2424 => x"83258403",
        2425 => x"63860500",
        2426 => x"13050400",
        2427 => x"ef000011",
        2428 => x"8325c403",
        2429 => x"63860500",
        2430 => x"13050400",
        2431 => x"ef000010",
        2432 => x"83250404",
        2433 => x"63860500",
        2434 => x"13050400",
        2435 => x"ef00000f",
        2436 => x"8325c405",
        2437 => x"63860500",
        2438 => x"13050400",
        2439 => x"ef00000e",
        2440 => x"83258405",
        2441 => x"63860500",
        2442 => x"13050400",
        2443 => x"ef00000d",
        2444 => x"83254403",
        2445 => x"63860500",
        2446 => x"13050400",
        2447 => x"ef00000c",
        2448 => x"83278401",
        2449 => x"638a0706",
        2450 => x"83278402",
        2451 => x"13050400",
        2452 => x"e7800700",
        2453 => x"83258404",
        2454 => x"63800506",
        2455 => x"13050400",
        2456 => x"03248101",
        2457 => x"8320c101",
        2458 => x"83244101",
        2459 => x"03290101",
        2460 => x"8329c100",
        2461 => x"13010102",
        2462 => x"6ff09feb",
        2463 => x"b3859500",
        2464 => x"83a50500",
        2465 => x"63900502",
        2466 => x"93844400",
        2467 => x"83274402",
        2468 => x"83a5c700",
        2469 => x"e39424ff",
        2470 => x"13050400",
        2471 => x"ef000006",
        2472 => x"6ff0dff0",
        2473 => x"83a90500",
        2474 => x"13050400",
        2475 => x"ef000005",
        2476 => x"93850900",
        2477 => x"6ff01ffd",
        2478 => x"8320c101",
        2479 => x"03248101",
        2480 => x"83244101",
        2481 => x"03290101",
        2482 => x"8329c100",
        2483 => x"13010102",
        2484 => x"67800000",
        2485 => x"67800000",
        2486 => x"93f5f50f",
        2487 => x"3306c500",
        2488 => x"6316c500",
        2489 => x"13050000",
        2490 => x"67800000",
        2491 => x"83470500",
        2492 => x"e38cb7fe",
        2493 => x"13051500",
        2494 => x"6ff09ffe",
        2495 => x"638a050e",
        2496 => x"83a7c5ff",
        2497 => x"130101fe",
        2498 => x"232c8100",
        2499 => x"232e1100",
        2500 => x"1384c5ff",
        2501 => x"63d40700",
        2502 => x"3304f400",
        2503 => x"2326a100",
        2504 => x"ef000034",
        2505 => x"83a78188",
        2506 => x"0325c100",
        2507 => x"639e0700",
        2508 => x"23220400",
        2509 => x"23a48188",
        2510 => x"03248101",
        2511 => x"8320c101",
        2512 => x"13010102",
        2513 => x"6f000032",
        2514 => x"6374f402",
        2515 => x"03260400",
        2516 => x"b306c400",
        2517 => x"639ad700",
        2518 => x"83a60700",
        2519 => x"83a74700",
        2520 => x"b386c600",
        2521 => x"2320d400",
        2522 => x"2322f400",
        2523 => x"6ff09ffc",
        2524 => x"13870700",
        2525 => x"83a74700",
        2526 => x"63840700",
        2527 => x"e37af4fe",
        2528 => x"83260700",
        2529 => x"3306d700",
        2530 => x"63188602",
        2531 => x"03260400",
        2532 => x"b386c600",
        2533 => x"2320d700",
        2534 => x"3306d700",
        2535 => x"e39ec7f8",
        2536 => x"03a60700",
        2537 => x"83a74700",
        2538 => x"b306d600",
        2539 => x"2320d700",
        2540 => x"2322f700",
        2541 => x"6ff05ff8",
        2542 => x"6378c400",
        2543 => x"9307c000",
        2544 => x"2320f500",
        2545 => x"6ff05ff7",
        2546 => x"03260400",
        2547 => x"b306c400",
        2548 => x"639ad700",
        2549 => x"83a60700",
        2550 => x"83a74700",
        2551 => x"b386c600",
        2552 => x"2320d400",
        2553 => x"2322f400",
        2554 => x"23228700",
        2555 => x"6ff0dff4",
        2556 => x"67800000",
        2557 => x"130101fe",
        2558 => x"232a9100",
        2559 => x"93843500",
        2560 => x"93f4c4ff",
        2561 => x"23282101",
        2562 => x"232e1100",
        2563 => x"232c8100",
        2564 => x"23263101",
        2565 => x"93848400",
        2566 => x"9307c000",
        2567 => x"13090500",
        2568 => x"63f4f406",
        2569 => x"9304c000",
        2570 => x"63e2b406",
        2571 => x"13050900",
        2572 => x"ef000023",
        2573 => x"03a78188",
        2574 => x"93868188",
        2575 => x"13040700",
        2576 => x"631a0406",
        2577 => x"1384c188",
        2578 => x"83270400",
        2579 => x"639a0700",
        2580 => x"93050000",
        2581 => x"13050900",
        2582 => x"ef00001c",
        2583 => x"2320a400",
        2584 => x"93850400",
        2585 => x"13050900",
        2586 => x"ef00001b",
        2587 => x"9309f0ff",
        2588 => x"631a350b",
        2589 => x"9307c000",
        2590 => x"2320f900",
        2591 => x"13050900",
        2592 => x"ef00401e",
        2593 => x"6f000001",
        2594 => x"e3d004fa",
        2595 => x"9307c000",
        2596 => x"2320f900",
        2597 => x"13050000",
        2598 => x"8320c101",
        2599 => x"03248101",
        2600 => x"83244101",
        2601 => x"03290101",
        2602 => x"8329c100",
        2603 => x"13010102",
        2604 => x"67800000",
        2605 => x"83270400",
        2606 => x"b3879740",
        2607 => x"63ce0704",
        2608 => x"1306b000",
        2609 => x"637af600",
        2610 => x"2320f400",
        2611 => x"3304f400",
        2612 => x"23209400",
        2613 => x"6f000001",
        2614 => x"83274400",
        2615 => x"631a8702",
        2616 => x"23a0f600",
        2617 => x"13050900",
        2618 => x"ef00c017",
        2619 => x"1305b400",
        2620 => x"93074400",
        2621 => x"137585ff",
        2622 => x"3307f540",
        2623 => x"e30ef5f8",
        2624 => x"3304e400",
        2625 => x"b387a740",
        2626 => x"2320f400",
        2627 => x"6ff0dff8",
        2628 => x"2322f700",
        2629 => x"6ff01ffd",
        2630 => x"13070400",
        2631 => x"03244400",
        2632 => x"6ff01ff2",
        2633 => x"13043500",
        2634 => x"1374c4ff",
        2635 => x"e30285fa",
        2636 => x"b305a440",
        2637 => x"13050900",
        2638 => x"ef00000e",
        2639 => x"e31a35f9",
        2640 => x"6ff05ff3",
        2641 => x"130101fe",
        2642 => x"232c8100",
        2643 => x"232e1100",
        2644 => x"232a9100",
        2645 => x"23282101",
        2646 => x"23263101",
        2647 => x"23244101",
        2648 => x"13040600",
        2649 => x"63940502",
        2650 => x"03248101",
        2651 => x"8320c101",
        2652 => x"83244101",
        2653 => x"03290101",
        2654 => x"8329c100",
        2655 => x"032a8100",
        2656 => x"93050600",
        2657 => x"13010102",
        2658 => x"6ff0dfe6",
        2659 => x"63180602",
        2660 => x"eff0dfd6",
        2661 => x"93040000",
        2662 => x"8320c101",
        2663 => x"03248101",
        2664 => x"03290101",
        2665 => x"8329c100",
        2666 => x"032a8100",
        2667 => x"13850400",
        2668 => x"83244101",
        2669 => x"13010102",
        2670 => x"67800000",
        2671 => x"130a0500",
        2672 => x"13890500",
        2673 => x"ef00400a",
        2674 => x"93090500",
        2675 => x"63688500",
        2676 => x"93571500",
        2677 => x"93040900",
        2678 => x"e3e087fc",
        2679 => x"93050400",
        2680 => x"13050a00",
        2681 => x"eff01fe1",
        2682 => x"93040500",
        2683 => x"e30605fa",
        2684 => x"13060400",
        2685 => x"63f48900",
        2686 => x"13860900",
        2687 => x"93050900",
        2688 => x"13850400",
        2689 => x"efe05f9d",
        2690 => x"93050900",
        2691 => x"13050a00",
        2692 => x"eff0dfce",
        2693 => x"6ff05ff8",
        2694 => x"130101ff",
        2695 => x"23248100",
        2696 => x"23229100",
        2697 => x"13040500",
        2698 => x"13850500",
        2699 => x"23261100",
        2700 => x"23a20188",
        2701 => x"ef00000c",
        2702 => x"9307f0ff",
        2703 => x"6318f500",
        2704 => x"83a74188",
        2705 => x"63840700",
        2706 => x"2320f400",
        2707 => x"8320c100",
        2708 => x"03248100",
        2709 => x"83244100",
        2710 => x"13010101",
        2711 => x"67800000",
        2712 => x"67800000",
        2713 => x"67800000",
        2714 => x"83a7c5ff",
        2715 => x"1385c7ff",
        2716 => x"63d80700",
        2717 => x"b385a500",
        2718 => x"83a70500",
        2719 => x"3305f500",
        2720 => x"67800000",
        2721 => x"9308d005",
        2722 => x"73000000",
        2723 => x"63520502",
        2724 => x"130101ff",
        2725 => x"23248100",
        2726 => x"13040500",
        2727 => x"23261100",
        2728 => x"33048040",
        2729 => x"efe05fc6",
        2730 => x"23208500",
        2731 => x"6f000000",
        2732 => x"6f000000",
        2733 => x"130101ff",
        2734 => x"23261100",
        2735 => x"23248100",
        2736 => x"9308900a",
        2737 => x"73000000",
        2738 => x"13040500",
        2739 => x"635a0500",
        2740 => x"33048040",
        2741 => x"efe05fc3",
        2742 => x"23208500",
        2743 => x"1304f0ff",
        2744 => x"8320c100",
        2745 => x"13050400",
        2746 => x"03248100",
        2747 => x"13010101",
        2748 => x"67800000",
        2749 => x"83a70189",
        2750 => x"130101ff",
        2751 => x"23261100",
        2752 => x"93060500",
        2753 => x"13870189",
        2754 => x"639c0702",
        2755 => x"9308600d",
        2756 => x"13050000",
        2757 => x"73000000",
        2758 => x"9307f0ff",
        2759 => x"6310f502",
        2760 => x"efe09fbe",
        2761 => x"9307c000",
        2762 => x"2320f500",
        2763 => x"1305f0ff",
        2764 => x"8320c100",
        2765 => x"13010101",
        2766 => x"67800000",
        2767 => x"2320a700",
        2768 => x"83270700",
        2769 => x"9308600d",
        2770 => x"b386f600",
        2771 => x"13850600",
        2772 => x"73000000",
        2773 => x"e316d5fc",
        2774 => x"2320a700",
        2775 => x"13850700",
        2776 => x"6ff01ffd",
        2777 => x"10000000",
        2778 => x"00000000",
        2779 => x"037a5200",
        2780 => x"017c0101",
        2781 => x"1b0d0200",
        2782 => x"10000000",
        2783 => x"18000000",
        2784 => x"ccdbffff",
        2785 => x"78040000",
        2786 => x"00000000",
        2787 => x"10000000",
        2788 => x"00000000",
        2789 => x"037a5200",
        2790 => x"017c0101",
        2791 => x"1b0d0200",
        2792 => x"10000000",
        2793 => x"18000000",
        2794 => x"1ce0ffff",
        2795 => x"30040000",
        2796 => x"00000000",
        2797 => x"10000000",
        2798 => x"00000000",
        2799 => x"037a5200",
        2800 => x"017c0101",
        2801 => x"1b0d0200",
        2802 => x"10000000",
        2803 => x"18000000",
        2804 => x"24e4ffff",
        2805 => x"e4030000",
        2806 => x"00000000",
        2807 => x"2c020000",
        2808 => x"9c010000",
        2809 => x"9c010000",
        2810 => x"9c010000",
        2811 => x"9c010000",
        2812 => x"10020000",
        2813 => x"9c010000",
        2814 => x"d0010000",
        2815 => x"9c010000",
        2816 => x"9c010000",
        2817 => x"d0010000",
        2818 => x"9c010000",
        2819 => x"9c010000",
        2820 => x"9c010000",
        2821 => x"9c010000",
        2822 => x"9c010000",
        2823 => x"9c010000",
        2824 => x"9c010000",
        2825 => x"80010000",
        2826 => x"28040000",
        2827 => x"28040000",
        2828 => x"28040000",
        2829 => x"80040000",
        2830 => x"28040000",
        2831 => x"28040000",
        2832 => x"28040000",
        2833 => x"28040000",
        2834 => x"28040000",
        2835 => x"28040000",
        2836 => x"28040000",
        2837 => x"48040000",
        2838 => x"ec040000",
        2839 => x"b4040000",
        2840 => x"b4040000",
        2841 => x"b4040000",
        2842 => x"b4040000",
        2843 => x"e0040000",
        2844 => x"74050000",
        2845 => x"4c050000",
        2846 => x"b4040000",
        2847 => x"b4040000",
        2848 => x"b4040000",
        2849 => x"b4040000",
        2850 => x"b4040000",
        2851 => x"b4040000",
        2852 => x"b4040000",
        2853 => x"b4040000",
        2854 => x"b4040000",
        2855 => x"b4040000",
        2856 => x"b4040000",
        2857 => x"b4040000",
        2858 => x"b4040000",
        2859 => x"b4040000",
        2860 => x"cc040000",
        2861 => x"cc040000",
        2862 => x"b4040000",
        2863 => x"b4040000",
        2864 => x"b4040000",
        2865 => x"b4040000",
        2866 => x"b4040000",
        2867 => x"b4040000",
        2868 => x"b4040000",
        2869 => x"b4040000",
        2870 => x"b4040000",
        2871 => x"b4040000",
        2872 => x"b4040000",
        2873 => x"b4040000",
        2874 => x"e0040000",
        2875 => x"ec040000",
        2876 => x"04050000",
        2877 => x"34050000",
        2878 => x"b4040000",
        2879 => x"b4040000",
        2880 => x"b4040000",
        2881 => x"b4040000",
        2882 => x"b4040000",
        2883 => x"b4040000",
        2884 => x"1c050000",
        2885 => x"b4040000",
        2886 => x"b4040000",
        2887 => x"b4040000",
        2888 => x"b4040000",
        2889 => x"cc040000",
        2890 => x"cc040000",
        2891 => x"00010202",
        2892 => x"03030303",
        2893 => x"04040404",
        2894 => x"04040404",
        2895 => x"05050505",
        2896 => x"05050505",
        2897 => x"05050505",
        2898 => x"05050505",
        2899 => x"06060606",
        2900 => x"06060606",
        2901 => x"06060606",
        2902 => x"06060606",
        2903 => x"06060606",
        2904 => x"06060606",
        2905 => x"06060606",
        2906 => x"06060606",
        2907 => x"07070707",
        2908 => x"07070707",
        2909 => x"07070707",
        2910 => x"07070707",
        2911 => x"07070707",
        2912 => x"07070707",
        2913 => x"07070707",
        2914 => x"07070707",
        2915 => x"07070707",
        2916 => x"07070707",
        2917 => x"07070707",
        2918 => x"07070707",
        2919 => x"07070707",
        2920 => x"07070707",
        2921 => x"07070707",
        2922 => x"07070707",
        2923 => x"08080808",
        2924 => x"08080808",
        2925 => x"08080808",
        2926 => x"08080808",
        2927 => x"08080808",
        2928 => x"08080808",
        2929 => x"08080808",
        2930 => x"08080808",
        2931 => x"08080808",
        2932 => x"08080808",
        2933 => x"08080808",
        2934 => x"08080808",
        2935 => x"08080808",
        2936 => x"08080808",
        2937 => x"08080808",
        2938 => x"08080808",
        2939 => x"08080808",
        2940 => x"08080808",
        2941 => x"08080808",
        2942 => x"08080808",
        2943 => x"08080808",
        2944 => x"08080808",
        2945 => x"08080808",
        2946 => x"08080808",
        2947 => x"08080808",
        2948 => x"08080808",
        2949 => x"08080808",
        2950 => x"08080808",
        2951 => x"08080808",
        2952 => x"08080808",
        2953 => x"08080808",
        2954 => x"08080808",
        2955 => x"0d0a0d0a",
        2956 => x"44697370",
        2957 => x"6c617969",
        2958 => x"6e672074",
        2959 => x"68652074",
        2960 => x"696d6520",
        2961 => x"70617373",
        2962 => x"65642073",
        2963 => x"696e6365",
        2964 => x"20726573",
        2965 => x"65740d0a",
        2966 => x"0d0a0000",
        2967 => x"2530356c",
        2968 => x"643a2530",
        2969 => x"366c6420",
        2970 => x"20202530",
        2971 => x"326c643a",
        2972 => x"2530326c",
        2973 => x"643a2530",
        2974 => x"326c640d",
        2975 => x"00000000",
        2976 => x"696e7465",
        2977 => x"72727570",
        2978 => x"745f6469",
        2979 => x"72656374",
        2980 => x"00000000",
        2981 => x"52495343",
        2982 => x"2d562052",
        2983 => x"56333249",
        2984 => x"4d206261",
        2985 => x"7265206d",
        2986 => x"6574616c",
        2987 => x"2070726f",
        2988 => x"63657373",
        2989 => x"6f720000",
        2990 => x"54686520",
        2991 => x"48616775",
        2992 => x"6520556e",
        2993 => x"69766572",
        2994 => x"73697479",
        2995 => x"206f6620",
        2996 => x"4170706c",
        2997 => x"69656420",
        2998 => x"53636965",
        2999 => x"6e636573",
        3000 => x"00000000",
        3001 => x"44657061",
        3002 => x"72746d65",
        3003 => x"6e74206f",
        3004 => x"6620456c",
        3005 => x"65637472",
        3006 => x"6963616c",
        3007 => x"20456e67",
        3008 => x"696e6565",
        3009 => x"72696e67",
        3010 => x"00000000",
        3011 => x"4a2e452e",
        3012 => x"4a2e206f",
        3013 => x"70206465",
        3014 => x"6e204272",
        3015 => x"6f757700",
        3016 => x"3c627265",
        3017 => x"616b3e0d",
        3018 => x"0a000000",
        3019 => x"0d0a4542",
        3020 => x"5245414b",
        3021 => x"21206d69",
        3022 => x"70203d20",
        3023 => x"00000000",
        3024 => x"232d302b",
        3025 => x"20000000",
        3026 => x"686c4c00",
        3027 => x"65666745",
        3028 => x"46470000",
        3029 => x"30313233",
        3030 => x"34353637",
        3031 => x"38394142",
        3032 => x"43444546",
        3033 => x"00000000",
        3034 => x"30313233",
        3035 => x"34353637",
        3036 => x"38396162",
        3037 => x"63646566",
        3038 => x"00000000",
        3039 => x"28220000",
        3040 => x"48220000",
        3041 => x"f4210000",
        3042 => x"f4210000",
        3043 => x"f4210000",
        3044 => x"f4210000",
        3045 => x"48220000",
        3046 => x"f4210000",
        3047 => x"f4210000",
        3048 => x"f4210000",
        3049 => x"f4210000",
        3050 => x"34240000",
        3051 => x"a0220000",
        3052 => x"b0230000",
        3053 => x"f4210000",
        3054 => x"f4210000",
        3055 => x"7c240000",
        3056 => x"f4210000",
        3057 => x"a0220000",
        3058 => x"f4210000",
        3059 => x"f4210000",
        3060 => x"bc230000",
        3061 => x"18000020",
        3062 => x"802e0000",
        3063 => x"942e0000",
        3064 => x"b82e0000",
        3065 => x"e42e0000",
        3066 => x"0c2f0000",
        3067 => x"00000000",
        3068 => x"00000000",
        3069 => x"00000000",
        3070 => x"00000000",
        3071 => x"00000000",
        3072 => x"00000000",
        3073 => x"00000000",
        3074 => x"00000000",
        3075 => x"00000000",
        3076 => x"00000000",
        3077 => x"00000000",
        3078 => x"00000000",
        3079 => x"00000000",
        3080 => x"00000000",
        3081 => x"00000000",
        3082 => x"00000000",
        3083 => x"00000000",
        3084 => x"00000000",
        3085 => x"00000000",
        3086 => x"00000000",
        3087 => x"00000000",
        3088 => x"00000000",
        3089 => x"00000000",
        3090 => x"00000000",
        3091 => x"00000000",
        3092 => x"80000020",
        3093 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
