-- srec2vhdl table generator
-- for input file main.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"93828206",
           6 => x"73905230",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef105009",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"93858538",
          21 => x"13050500",
          22 => x"ef10d004",
          23 => x"ef10502b",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10100b",
          29 => x"ef10d025",
          30 => x"6f000000",
          31 => x"37170000",
          32 => x"b70700f0",
          33 => x"13077745",
          34 => x"23a2e702",
          35 => x"13070004",
          36 => x"23a4e702",
          37 => x"67800000",
          38 => x"1375f50f",
          39 => x"b70700f0",
          40 => x"23a0a702",
          41 => x"370700f0",
          42 => x"8327c702",
          43 => x"93f70701",
          44 => x"e38c07fe",
          45 => x"67800000",
          46 => x"63060502",
          47 => x"83470500",
          48 => x"63820702",
          49 => x"370700f0",
          50 => x"13051500",
          51 => x"2320f702",
          52 => x"8327c702",
          53 => x"93f70701",
          54 => x"e38c07fe",
          55 => x"83470500",
          56 => x"e39407fe",
          57 => x"67800000",
          58 => x"370700f0",
          59 => x"8327c702",
          60 => x"93f74700",
          61 => x"e38c07fe",
          62 => x"03250702",
          63 => x"1375f50f",
          64 => x"67800000",
          65 => x"130101ff",
          66 => x"373e0000",
          67 => x"370700f0",
          68 => x"930e0500",
          69 => x"138ff5ff",
          70 => x"23268100",
          71 => x"13050000",
          72 => x"130e4efc",
          73 => x"13070702",
          74 => x"13035001",
          75 => x"93027000",
          76 => x"930fe005",
          77 => x"9305f007",
          78 => x"93082000",
          79 => x"13082001",
          80 => x"b7330000",
          81 => x"1306f007",
          82 => x"8327c700",
          83 => x"93f74700",
          84 => x"e38c07fe",
          85 => x"03240700",
          86 => x"9376f40f",
          87 => x"636ed302",
          88 => x"63fed802",
          89 => x"9387d6ff",
          90 => x"636af802",
          91 => x"93972700",
          92 => x"b307fe00",
          93 => x"83a70700",
          94 => x"67800700",
          95 => x"1305f5ff",
          96 => x"6308050c",
          97 => x"2320c700",
          98 => x"8327c700",
          99 => x"93f70701",
         100 => x"e38c07fe",
         101 => x"6ff09ffe",
         102 => x"638cb606",
         103 => x"635ae50d",
         104 => x"1374f40f",
         105 => x"930704fe",
         106 => x"93f7f70f",
         107 => x"e3eefff8",
         108 => x"b387ae00",
         109 => x"23808700",
         110 => x"13051500",
         111 => x"2320d700",
         112 => x"8327c700",
         113 => x"93f70701",
         114 => x"e38c07fe",
         115 => x"6ff0dff7",
         116 => x"b38eae00",
         117 => x"b7360000",
         118 => x"23800e00",
         119 => x"9307d000",
         120 => x"93860621",
         121 => x"370700f0",
         122 => x"93861600",
         123 => x"2320f702",
         124 => x"8327c702",
         125 => x"93f70701",
         126 => x"e38c07fe",
         127 => x"83c70600",
         128 => x"e39407fe",
         129 => x"0324c100",
         130 => x"13010101",
         131 => x"67800000",
         132 => x"63040504",
         133 => x"2320b700",
         134 => x"8327c700",
         135 => x"93f70701",
         136 => x"e38c07fe",
         137 => x"1305f5ff",
         138 => x"6ff01ff2",
         139 => x"9307c003",
         140 => x"9386032d",
         141 => x"93861600",
         142 => x"2320f700",
         143 => x"8327c700",
         144 => x"93f70701",
         145 => x"e38c07fe",
         146 => x"83c70600",
         147 => x"e39407fe",
         148 => x"13050000",
         149 => x"6ff05fef",
         150 => x"23205700",
         151 => x"8327c700",
         152 => x"93f70701",
         153 => x"e38c07fe",
         154 => x"13050000",
         155 => x"6ff0dfed",
         156 => x"23205700",
         157 => x"8327c700",
         158 => x"93f70701",
         159 => x"e38c07fe",
         160 => x"6ff09fec",
         161 => x"1375f50f",
         162 => x"b70700f0",
         163 => x"23a0a702",
         164 => x"370700f0",
         165 => x"8327c702",
         166 => x"93f70701",
         167 => x"e38c07fe",
         168 => x"13051000",
         169 => x"67800000",
         170 => x"370700f0",
         171 => x"8327c702",
         172 => x"93f74700",
         173 => x"e38c07fe",
         174 => x"03250702",
         175 => x"1375f50f",
         176 => x"67800000",
         177 => x"13050000",
         178 => x"67800000",
         179 => x"13050000",
         180 => x"67800000",
         181 => x"6f000008",
         182 => x"6f004043",
         183 => x"6f000043",
         184 => x"6f00c042",
         185 => x"6f008042",
         186 => x"6f004042",
         187 => x"6f000042",
         188 => x"6f000042",
         189 => x"6f008041",
         190 => x"6f004041",
         191 => x"6f000041",
         192 => x"6f00c040",
         193 => x"6f008040",
         194 => x"6f004040",
         195 => x"6f000040",
         196 => x"6f00c03f",
         197 => x"6f00803f",
         198 => x"6f00403b",
         199 => x"6f000047",
         200 => x"6f00c03e",
         201 => x"6f00803e",
         202 => x"6f00403e",
         203 => x"6f00003e",
         204 => x"6f00c03d",
         205 => x"6f00803d",
         206 => x"6f00403d",
         207 => x"6f00003d",
         208 => x"6f00c03c",
         209 => x"6f00803c",
         210 => x"6f00403c",
         211 => x"6f00003c",
         212 => x"6f00c03b",
         213 => x"130101f8",
         214 => x"23221100",
         215 => x"23242100",
         216 => x"23263100",
         217 => x"23284100",
         218 => x"232a5100",
         219 => x"232c6100",
         220 => x"232e7100",
         221 => x"23208102",
         222 => x"23229102",
         223 => x"2324a102",
         224 => x"2326b102",
         225 => x"2328c102",
         226 => x"232ad102",
         227 => x"232ce102",
         228 => x"232ef102",
         229 => x"23200105",
         230 => x"23221105",
         231 => x"23242105",
         232 => x"23263105",
         233 => x"23284105",
         234 => x"232a5105",
         235 => x"232c6105",
         236 => x"232e7105",
         237 => x"23208107",
         238 => x"23229107",
         239 => x"2324a107",
         240 => x"2326b107",
         241 => x"2328c107",
         242 => x"232ad107",
         243 => x"232ce107",
         244 => x"232ef107",
         245 => x"f3272034",
         246 => x"1307b000",
         247 => x"6388e708",
         248 => x"13073000",
         249 => x"638ce70e",
         250 => x"03258102",
         251 => x"832fc107",
         252 => x"032f8107",
         253 => x"832e4107",
         254 => x"032e0107",
         255 => x"832dc106",
         256 => x"032d8106",
         257 => x"832c4106",
         258 => x"032c0106",
         259 => x"832bc105",
         260 => x"032b8105",
         261 => x"832a4105",
         262 => x"032a0105",
         263 => x"8329c104",
         264 => x"03298104",
         265 => x"83284104",
         266 => x"03280104",
         267 => x"8327c103",
         268 => x"03278103",
         269 => x"83264103",
         270 => x"03260103",
         271 => x"8325c102",
         272 => x"83244102",
         273 => x"03240102",
         274 => x"8323c101",
         275 => x"03238101",
         276 => x"83224101",
         277 => x"03220101",
         278 => x"8321c100",
         279 => x"03218100",
         280 => x"83204100",
         281 => x"13010108",
         282 => x"73002030",
         283 => x"9307600d",
         284 => x"638ef806",
         285 => x"9307900a",
         286 => x"6382f818",
         287 => x"63c41703",
         288 => x"938878fc",
         289 => x"93074002",
         290 => x"63e0170b",
         291 => x"b7370000",
         292 => x"93870701",
         293 => x"93982800",
         294 => x"b388f800",
         295 => x"83a70800",
         296 => x"67800700",
         297 => x"938808c0",
         298 => x"9307f000",
         299 => x"63ee1707",
         300 => x"b7370000",
         301 => x"9387470a",
         302 => x"93982800",
         303 => x"b388f800",
         304 => x"83a70800",
         305 => x"67800700",
         306 => x"b7270000",
         307 => x"23a2f500",
         308 => x"93070000",
         309 => x"13850700",
         310 => x"6ff05ff1",
         311 => x"13050100",
         312 => x"ef004018",
         313 => x"03258102",
         314 => x"6ff05ff0",
         315 => x"63180500",
         316 => x"13858189",
         317 => x"13050500",
         318 => x"6ff05fef",
         319 => x"b7870020",
         320 => x"93870700",
         321 => x"13070040",
         322 => x"b387e740",
         323 => x"e364f5fe",
         324 => x"ef10805b",
         325 => x"9307c000",
         326 => x"2320f500",
         327 => x"1305f0ff",
         328 => x"13050500",
         329 => x"6ff09fec",
         330 => x"ef10005a",
         331 => x"93078005",
         332 => x"2320f500",
         333 => x"9307f0ff",
         334 => x"13850700",
         335 => x"6ff01feb",
         336 => x"ef108058",
         337 => x"93079000",
         338 => x"2320f500",
         339 => x"9307f0ff",
         340 => x"13850700",
         341 => x"6ff09fe9",
         342 => x"93070000",
         343 => x"13850700",
         344 => x"6ff0dfe8",
         345 => x"ef104056",
         346 => x"9307d000",
         347 => x"2320f500",
         348 => x"9307f0ff",
         349 => x"13850700",
         350 => x"6ff05fe7",
         351 => x"ef10c054",
         352 => x"9307f001",
         353 => x"2320f500",
         354 => x"9307f0ff",
         355 => x"13850700",
         356 => x"6ff0dfe5",
         357 => x"ef104053",
         358 => x"93072000",
         359 => x"2320f500",
         360 => x"9307f0ff",
         361 => x"13850700",
         362 => x"6ff05fe4",
         363 => x"13090600",
         364 => x"13840500",
         365 => x"635cc000",
         366 => x"b384c500",
         367 => x"eff0dfce",
         368 => x"2300a400",
         369 => x"13041400",
         370 => x"e31a94fe",
         371 => x"13050900",
         372 => x"6ff0dfe1",
         373 => x"13090600",
         374 => x"13840500",
         375 => x"e358c0fe",
         376 => x"b384c500",
         377 => x"03450400",
         378 => x"13041400",
         379 => x"eff09fc9",
         380 => x"e39a84fe",
         381 => x"13050900",
         382 => x"6ff05fdf",
         383 => x"13090000",
         384 => x"93040500",
         385 => x"13040900",
         386 => x"93090900",
         387 => x"93070900",
         388 => x"732410c8",
         389 => x"f32910c0",
         390 => x"f32710c8",
         391 => x"e31af4fe",
         392 => x"37460f00",
         393 => x"13060624",
         394 => x"93060000",
         395 => x"13850900",
         396 => x"93050400",
         397 => x"ef00d068",
         398 => x"37460f00",
         399 => x"23a4a400",
         400 => x"13060624",
         401 => x"93060000",
         402 => x"13850900",
         403 => x"93050400",
         404 => x"ef001024",
         405 => x"23a0a400",
         406 => x"23a2b400",
         407 => x"13050900",
         408 => x"6ff0dfd8",
         409 => x"37350000",
         410 => x"130101ff",
         411 => x"1305c52d",
         412 => x"23261100",
         413 => x"23248100",
         414 => x"23229100",
         415 => x"23202101",
         416 => x"eff09fa3",
         417 => x"73294034",
         418 => x"93040002",
         419 => x"37040080",
         420 => x"33758900",
         421 => x"3335a000",
         422 => x"13050503",
         423 => x"9384f4ff",
         424 => x"eff09f9f",
         425 => x"13541400",
         426 => x"e39404fe",
         427 => x"03248100",
         428 => x"8320c100",
         429 => x"83244100",
         430 => x"03290100",
         431 => x"37350000",
         432 => x"13050521",
         433 => x"13010101",
         434 => x"6ff01f9f",
         435 => x"130101ff",
         436 => x"2322f100",
         437 => x"b70700f0",
         438 => x"2324e100",
         439 => x"03a74708",
         440 => x"2326d100",
         441 => x"8326c100",
         442 => x"1377f7fe",
         443 => x"23a2e708",
         444 => x"03a74700",
         445 => x"13471700",
         446 => x"23a2e700",
         447 => x"03278100",
         448 => x"83274100",
         449 => x"13010101",
         450 => x"73002030",
         451 => x"6f000000",
         452 => x"130101fe",
         453 => x"2326f100",
         454 => x"232eb100",
         455 => x"232cc100",
         456 => x"232ad100",
         457 => x"2328e100",
         458 => x"b70700f0",
         459 => x"83a6470f",
         460 => x"03a6070f",
         461 => x"03a7470f",
         462 => x"e31ad7fe",
         463 => x"b7860100",
         464 => x"9305f0ff",
         465 => x"9386066a",
         466 => x"23aeb70e",
         467 => x"b306d600",
         468 => x"23acb70e",
         469 => x"33b6c600",
         470 => x"23acd70e",
         471 => x"3306e600",
         472 => x"23aec70e",
         473 => x"03a74700",
         474 => x"8325c101",
         475 => x"03268101",
         476 => x"13472700",
         477 => x"23a2e700",
         478 => x"83264101",
         479 => x"03270101",
         480 => x"8327c100",
         481 => x"13010102",
         482 => x"73002030",
         483 => x"130101ff",
         484 => x"2326e100",
         485 => x"370700f0",
         486 => x"2324f100",
         487 => x"8327c702",
         488 => x"93f74700",
         489 => x"638a0700",
         490 => x"83274700",
         491 => x"93c74700",
         492 => x"2322f700",
         493 => x"83270702",
         494 => x"0327c100",
         495 => x"83278100",
         496 => x"13010101",
         497 => x"73002030",
         498 => x"13030500",
         499 => x"138e0500",
         500 => x"93080000",
         501 => x"63dc0500",
         502 => x"b337a000",
         503 => x"330eb040",
         504 => x"330efe40",
         505 => x"3303a040",
         506 => x"9308f0ff",
         507 => x"63dc0600",
         508 => x"b337c000",
         509 => x"b306d040",
         510 => x"93c8f8ff",
         511 => x"b386f640",
         512 => x"3306c040",
         513 => x"13070600",
         514 => x"13080300",
         515 => x"93070e00",
         516 => x"639c0628",
         517 => x"b7350000",
         518 => x"9385450e",
         519 => x"6376ce0e",
         520 => x"b7060100",
         521 => x"6378d60c",
         522 => x"93360610",
         523 => x"93c61600",
         524 => x"93963600",
         525 => x"3355d600",
         526 => x"b385a500",
         527 => x"83c50500",
         528 => x"13050002",
         529 => x"b386d500",
         530 => x"b305d540",
         531 => x"630cd500",
         532 => x"b317be00",
         533 => x"b356d300",
         534 => x"3317b600",
         535 => x"b3e7f600",
         536 => x"3318b300",
         537 => x"93550701",
         538 => x"33deb702",
         539 => x"13160701",
         540 => x"13560601",
         541 => x"b3f7b702",
         542 => x"13050e00",
         543 => x"3303c603",
         544 => x"93960701",
         545 => x"93570801",
         546 => x"b3e7d700",
         547 => x"63fe6700",
         548 => x"b387e700",
         549 => x"1305feff",
         550 => x"63e8e700",
         551 => x"63f66700",
         552 => x"1305eeff",
         553 => x"b387e700",
         554 => x"b3876740",
         555 => x"33d3b702",
         556 => x"13180801",
         557 => x"13580801",
         558 => x"b3f7b702",
         559 => x"b3066602",
         560 => x"93970701",
         561 => x"3368f800",
         562 => x"93070300",
         563 => x"637cd800",
         564 => x"33080701",
         565 => x"9307f3ff",
         566 => x"6366e800",
         567 => x"6374d800",
         568 => x"9307e3ff",
         569 => x"13150501",
         570 => x"3365f500",
         571 => x"93050000",
         572 => x"6f00000e",
         573 => x"37050001",
         574 => x"93060001",
         575 => x"e36ca6f2",
         576 => x"93068001",
         577 => x"6ff01ff3",
         578 => x"63140600",
         579 => x"73001000",
         580 => x"b7070100",
         581 => x"637af60c",
         582 => x"93360610",
         583 => x"93c61600",
         584 => x"93963600",
         585 => x"b357d600",
         586 => x"b385f500",
         587 => x"83c70500",
         588 => x"b387d700",
         589 => x"93060002",
         590 => x"b385f640",
         591 => x"6390f60c",
         592 => x"b307ce40",
         593 => x"93051000",
         594 => x"13530701",
         595 => x"b3de6702",
         596 => x"13160701",
         597 => x"13560601",
         598 => x"93560801",
         599 => x"b3f76702",
         600 => x"13850e00",
         601 => x"330ed603",
         602 => x"93970701",
         603 => x"b3e7f600",
         604 => x"63fec701",
         605 => x"b387e700",
         606 => x"1385feff",
         607 => x"63e8e700",
         608 => x"63f6c701",
         609 => x"1385eeff",
         610 => x"b387e700",
         611 => x"b387c741",
         612 => x"33de6702",
         613 => x"13180801",
         614 => x"13580801",
         615 => x"b3f76702",
         616 => x"b306c603",
         617 => x"93970701",
         618 => x"3368f800",
         619 => x"93070e00",
         620 => x"637cd800",
         621 => x"33080701",
         622 => x"9307feff",
         623 => x"6366e800",
         624 => x"6374d800",
         625 => x"9307eeff",
         626 => x"13150501",
         627 => x"3365f500",
         628 => x"638a0800",
         629 => x"b337a000",
         630 => x"b305b040",
         631 => x"b385f540",
         632 => x"3305a040",
         633 => x"67800000",
         634 => x"b7070001",
         635 => x"93060001",
         636 => x"e36af6f2",
         637 => x"93068001",
         638 => x"6ff0dff2",
         639 => x"3317b600",
         640 => x"b356fe00",
         641 => x"13550701",
         642 => x"331ebe00",
         643 => x"b357f300",
         644 => x"b3e7c701",
         645 => x"33dea602",
         646 => x"13160701",
         647 => x"13560601",
         648 => x"3318b300",
         649 => x"b3f6a602",
         650 => x"3303c603",
         651 => x"93950601",
         652 => x"93d60701",
         653 => x"b3e6b600",
         654 => x"93050e00",
         655 => x"63fe6600",
         656 => x"b386e600",
         657 => x"9305feff",
         658 => x"63e8e600",
         659 => x"63f66600",
         660 => x"9305eeff",
         661 => x"b386e600",
         662 => x"b3866640",
         663 => x"33d3a602",
         664 => x"93970701",
         665 => x"93d70701",
         666 => x"b3f6a602",
         667 => x"33066602",
         668 => x"93960601",
         669 => x"b3e7d700",
         670 => x"93060300",
         671 => x"63fec700",
         672 => x"b387e700",
         673 => x"9306f3ff",
         674 => x"63e8e700",
         675 => x"63f6c700",
         676 => x"9306e3ff",
         677 => x"b387e700",
         678 => x"93950501",
         679 => x"b387c740",
         680 => x"b3e5d500",
         681 => x"6ff05fea",
         682 => x"6366de18",
         683 => x"b7070100",
         684 => x"63f4f604",
         685 => x"13b70610",
         686 => x"13471700",
         687 => x"13173700",
         688 => x"b7370000",
         689 => x"b3d5e600",
         690 => x"9387470e",
         691 => x"b387b700",
         692 => x"83c70700",
         693 => x"b387e700",
         694 => x"13070002",
         695 => x"b305f740",
         696 => x"6316f702",
         697 => x"13051000",
         698 => x"e3e4c6ef",
         699 => x"3335c300",
         700 => x"13451500",
         701 => x"6ff0dfed",
         702 => x"b7070001",
         703 => x"13070001",
         704 => x"e3e0f6fc",
         705 => x"13078001",
         706 => x"6ff09ffb",
         707 => x"3357f600",
         708 => x"b396b600",
         709 => x"b366d700",
         710 => x"3357fe00",
         711 => x"331ebe00",
         712 => x"b357f300",
         713 => x"b3e7c701",
         714 => x"13de0601",
         715 => x"335fc703",
         716 => x"13980601",
         717 => x"13580801",
         718 => x"3316b600",
         719 => x"3377c703",
         720 => x"b30ee803",
         721 => x"13150701",
         722 => x"13d70701",
         723 => x"3367a700",
         724 => x"13050f00",
         725 => x"637ed701",
         726 => x"3307d700",
         727 => x"1305ffff",
         728 => x"6368d700",
         729 => x"6376d701",
         730 => x"1305efff",
         731 => x"3307d700",
         732 => x"3307d741",
         733 => x"b35ec703",
         734 => x"93970701",
         735 => x"93d70701",
         736 => x"3377c703",
         737 => x"3308d803",
         738 => x"13170701",
         739 => x"b3e7e700",
         740 => x"13870e00",
         741 => x"63fe0701",
         742 => x"b387d700",
         743 => x"1387feff",
         744 => x"63e8d700",
         745 => x"63f60701",
         746 => x"1387eeff",
         747 => x"b387d700",
         748 => x"13150501",
         749 => x"b70e0100",
         750 => x"3365e500",
         751 => x"9386feff",
         752 => x"3377d500",
         753 => x"b3870741",
         754 => x"b376d600",
         755 => x"13580501",
         756 => x"13560601",
         757 => x"330ed702",
         758 => x"b306d802",
         759 => x"3307c702",
         760 => x"3308c802",
         761 => x"3306d700",
         762 => x"13570e01",
         763 => x"3307c700",
         764 => x"6374d700",
         765 => x"3308d801",
         766 => x"93560701",
         767 => x"b3860601",
         768 => x"63e6d702",
         769 => x"e394d7ce",
         770 => x"b7070100",
         771 => x"9387f7ff",
         772 => x"3377f700",
         773 => x"13170701",
         774 => x"337efe00",
         775 => x"3313b300",
         776 => x"3307c701",
         777 => x"93050000",
         778 => x"e374e3da",
         779 => x"1305f5ff",
         780 => x"6ff0dfcb",
         781 => x"93050000",
         782 => x"13050000",
         783 => x"6ff05fd9",
         784 => x"138e0500",
         785 => x"13080000",
         786 => x"63dc0500",
         787 => x"b337a000",
         788 => x"b305b040",
         789 => x"338ef540",
         790 => x"3305a040",
         791 => x"1308f0ff",
         792 => x"63da0600",
         793 => x"b337c000",
         794 => x"b306d040",
         795 => x"b386f640",
         796 => x"3306c040",
         797 => x"93080600",
         798 => x"93070500",
         799 => x"93050e00",
         800 => x"63940624",
         801 => x"37370000",
         802 => x"1307470e",
         803 => x"6376ce0e",
         804 => x"b7060100",
         805 => x"6378d60c",
         806 => x"93360610",
         807 => x"93c61600",
         808 => x"93963600",
         809 => x"3353d600",
         810 => x"33076700",
         811 => x"03470700",
         812 => x"3307d700",
         813 => x"93060002",
         814 => x"3383e640",
         815 => x"638ce600",
         816 => x"b3156e00",
         817 => x"3357e500",
         818 => x"b3186600",
         819 => x"b365b700",
         820 => x"b3176500",
         821 => x"93d60801",
         822 => x"33d7d502",
         823 => x"13950801",
         824 => x"13550501",
         825 => x"b3f5d502",
         826 => x"3307a702",
         827 => x"13960501",
         828 => x"93d50701",
         829 => x"b3e5c500",
         830 => x"63fae500",
         831 => x"b3851501",
         832 => x"63e61501",
         833 => x"63f4e500",
         834 => x"b3851501",
         835 => x"b385e540",
         836 => x"33d7d502",
         837 => x"93970701",
         838 => x"93d70701",
         839 => x"b3f5d502",
         840 => x"3307a702",
         841 => x"93950501",
         842 => x"b3e7b700",
         843 => x"63fae700",
         844 => x"b3871701",
         845 => x"63e61701",
         846 => x"63f4e700",
         847 => x"b3871701",
         848 => x"b387e740",
         849 => x"33d56700",
         850 => x"93050000",
         851 => x"630a0800",
         852 => x"b337a000",
         853 => x"b305b040",
         854 => x"b385f540",
         855 => x"3305a040",
         856 => x"67800000",
         857 => x"37030001",
         858 => x"93060001",
         859 => x"e36c66f2",
         860 => x"93068001",
         861 => x"6ff01ff3",
         862 => x"63140600",
         863 => x"73001000",
         864 => x"b7060100",
         865 => x"6372d60a",
         866 => x"93360610",
         867 => x"93c61600",
         868 => x"93963600",
         869 => x"b355d600",
         870 => x"3307b700",
         871 => x"03470700",
         872 => x"3307d700",
         873 => x"93060002",
         874 => x"3383e640",
         875 => x"6398e608",
         876 => x"3307ce40",
         877 => x"93d50801",
         878 => x"3356b702",
         879 => x"13950801",
         880 => x"13550501",
         881 => x"93d60701",
         882 => x"3377b702",
         883 => x"3306a602",
         884 => x"13170701",
         885 => x"33e7e600",
         886 => x"637ac700",
         887 => x"33071701",
         888 => x"63661701",
         889 => x"6374c700",
         890 => x"33071701",
         891 => x"3307c740",
         892 => x"b356b702",
         893 => x"93970701",
         894 => x"93d70701",
         895 => x"3377b702",
         896 => x"b386a602",
         897 => x"13170701",
         898 => x"b3e7e700",
         899 => x"63fad700",
         900 => x"b3871701",
         901 => x"63e61701",
         902 => x"63f4d700",
         903 => x"b3871701",
         904 => x"b387d740",
         905 => x"6ff01ff2",
         906 => x"b7050001",
         907 => x"93060001",
         908 => x"e362b6f6",
         909 => x"93068001",
         910 => x"6ff0dff5",
         911 => x"b3186600",
         912 => x"b356ee00",
         913 => x"b3156e00",
         914 => x"3357e500",
         915 => x"b3176500",
         916 => x"13d50801",
         917 => x"3367b700",
         918 => x"b3d5a602",
         919 => x"139e0801",
         920 => x"135e0e01",
         921 => x"b3f6a602",
         922 => x"b385c503",
         923 => x"13960601",
         924 => x"93560701",
         925 => x"b3e6c600",
         926 => x"63fab600",
         927 => x"b3861601",
         928 => x"63e61601",
         929 => x"63f4b600",
         930 => x"b3861601",
         931 => x"b386b640",
         932 => x"33d6a602",
         933 => x"13170701",
         934 => x"13570701",
         935 => x"b3f6a602",
         936 => x"3306c603",
         937 => x"93960601",
         938 => x"3367d700",
         939 => x"637ac700",
         940 => x"33071701",
         941 => x"63661701",
         942 => x"6374c700",
         943 => x"33071701",
         944 => x"3307c740",
         945 => x"6ff01fef",
         946 => x"e362dee8",
         947 => x"37070100",
         948 => x"63fce604",
         949 => x"13b70610",
         950 => x"13471700",
         951 => x"13173700",
         952 => x"b7380000",
         953 => x"33d3e600",
         954 => x"9388480e",
         955 => x"b3886800",
         956 => x"03c30800",
         957 => x"3303e300",
         958 => x"13070002",
         959 => x"b3086740",
         960 => x"631e6702",
         961 => x"63e4c601",
         962 => x"636cc500",
         963 => x"3306c540",
         964 => x"b306de40",
         965 => x"b335c500",
         966 => x"b385b640",
         967 => x"93070600",
         968 => x"13850700",
         969 => x"6ff09fe2",
         970 => x"b7080001",
         971 => x"13070001",
         972 => x"e3e816fb",
         973 => x"13078001",
         974 => x"6ff09ffa",
         975 => x"b3576600",
         976 => x"b3961601",
         977 => x"b3e6d700",
         978 => x"33576e00",
         979 => x"93de0601",
         980 => x"b35fd703",
         981 => x"b3151e01",
         982 => x"139e0601",
         983 => x"135e0e01",
         984 => x"b3576500",
         985 => x"b3e5b700",
         986 => x"93d70501",
         987 => x"33161601",
         988 => x"33151501",
         989 => x"3377d703",
         990 => x"330ffe03",
         991 => x"13170701",
         992 => x"b3e7e700",
         993 => x"13870f00",
         994 => x"63fee701",
         995 => x"b387d700",
         996 => x"1387ffff",
         997 => x"63e8d700",
         998 => x"63f6e701",
         999 => x"1387efff",
        1000 => x"b387d700",
        1001 => x"b387e741",
        1002 => x"33dfd703",
        1003 => x"93950501",
        1004 => x"93d50501",
        1005 => x"b3f7d703",
        1006 => x"330eee03",
        1007 => x"93970701",
        1008 => x"b3e5f500",
        1009 => x"93070f00",
        1010 => x"63fec501",
        1011 => x"b385d500",
        1012 => x"9307ffff",
        1013 => x"63e8d500",
        1014 => x"63f6c501",
        1015 => x"9307efff",
        1016 => x"b385d500",
        1017 => x"13170701",
        1018 => x"b70f0100",
        1019 => x"3367f700",
        1020 => x"b385c541",
        1021 => x"138effff",
        1022 => x"b377c701",
        1023 => x"935e0601",
        1024 => x"13570701",
        1025 => x"337ec601",
        1026 => x"338fc703",
        1027 => x"330ec703",
        1028 => x"b387d703",
        1029 => x"3307d703",
        1030 => x"b38ec701",
        1031 => x"93570f01",
        1032 => x"b387d701",
        1033 => x"63f4c701",
        1034 => x"3307f701",
        1035 => x"13de0701",
        1036 => x"3307ee00",
        1037 => x"370e0100",
        1038 => x"130efeff",
        1039 => x"b3f7c701",
        1040 => x"93970701",
        1041 => x"337fcf01",
        1042 => x"b387e701",
        1043 => x"63e6e500",
        1044 => x"639ee500",
        1045 => x"637cf500",
        1046 => x"3386c740",
        1047 => x"b3b7c700",
        1048 => x"b387d700",
        1049 => x"3307f740",
        1050 => x"93070600",
        1051 => x"b307f540",
        1052 => x"3335f500",
        1053 => x"b385e540",
        1054 => x"b385a540",
        1055 => x"33936500",
        1056 => x"b3d71701",
        1057 => x"3365f300",
        1058 => x"b3d51501",
        1059 => x"6ff01fcc",
        1060 => x"13030500",
        1061 => x"93880500",
        1062 => x"13070600",
        1063 => x"13080500",
        1064 => x"93870500",
        1065 => x"63920628",
        1066 => x"b7350000",
        1067 => x"9385450e",
        1068 => x"63f6c80e",
        1069 => x"b7060100",
        1070 => x"6378d60c",
        1071 => x"93360610",
        1072 => x"93c61600",
        1073 => x"93963600",
        1074 => x"3355d600",
        1075 => x"b385a500",
        1076 => x"83c50500",
        1077 => x"13050002",
        1078 => x"b386d500",
        1079 => x"b305d540",
        1080 => x"630cd500",
        1081 => x"b397b800",
        1082 => x"b356d300",
        1083 => x"3317b600",
        1084 => x"b3e7f600",
        1085 => x"3318b300",
        1086 => x"93550701",
        1087 => x"33d3b702",
        1088 => x"13160701",
        1089 => x"13560601",
        1090 => x"b3f7b702",
        1091 => x"13050300",
        1092 => x"b3086602",
        1093 => x"93960701",
        1094 => x"93570801",
        1095 => x"b3e7d700",
        1096 => x"63fe1701",
        1097 => x"b387e700",
        1098 => x"1305f3ff",
        1099 => x"63e8e700",
        1100 => x"63f61701",
        1101 => x"1305e3ff",
        1102 => x"b387e700",
        1103 => x"b3871741",
        1104 => x"b3d8b702",
        1105 => x"13180801",
        1106 => x"13580801",
        1107 => x"b3f7b702",
        1108 => x"b3061603",
        1109 => x"93970701",
        1110 => x"3368f800",
        1111 => x"93870800",
        1112 => x"637cd800",
        1113 => x"33080701",
        1114 => x"9387f8ff",
        1115 => x"6366e800",
        1116 => x"6374d800",
        1117 => x"9387e8ff",
        1118 => x"13150501",
        1119 => x"3365f500",
        1120 => x"93050000",
        1121 => x"67800000",
        1122 => x"37050001",
        1123 => x"93060001",
        1124 => x"e36ca6f2",
        1125 => x"93068001",
        1126 => x"6ff01ff3",
        1127 => x"63140600",
        1128 => x"73001000",
        1129 => x"b7070100",
        1130 => x"6370f60c",
        1131 => x"93360610",
        1132 => x"93c61600",
        1133 => x"93963600",
        1134 => x"b357d600",
        1135 => x"b385f500",
        1136 => x"83c70500",
        1137 => x"b387d700",
        1138 => x"93060002",
        1139 => x"b385f640",
        1140 => x"6396f60a",
        1141 => x"b387c840",
        1142 => x"93051000",
        1143 => x"93580701",
        1144 => x"33de1703",
        1145 => x"13160701",
        1146 => x"13560601",
        1147 => x"93560801",
        1148 => x"b3f71703",
        1149 => x"13050e00",
        1150 => x"3303c603",
        1151 => x"93970701",
        1152 => x"b3e7f600",
        1153 => x"63fe6700",
        1154 => x"b387e700",
        1155 => x"1305feff",
        1156 => x"63e8e700",
        1157 => x"63f66700",
        1158 => x"1305eeff",
        1159 => x"b387e700",
        1160 => x"b3876740",
        1161 => x"33d31703",
        1162 => x"13180801",
        1163 => x"13580801",
        1164 => x"b3f71703",
        1165 => x"b3066602",
        1166 => x"93970701",
        1167 => x"3368f800",
        1168 => x"93070300",
        1169 => x"637cd800",
        1170 => x"33080701",
        1171 => x"9307f3ff",
        1172 => x"6366e800",
        1173 => x"6374d800",
        1174 => x"9307e3ff",
        1175 => x"13150501",
        1176 => x"3365f500",
        1177 => x"67800000",
        1178 => x"b7070001",
        1179 => x"93060001",
        1180 => x"e364f6f4",
        1181 => x"93068001",
        1182 => x"6ff01ff4",
        1183 => x"3317b600",
        1184 => x"b3d6f800",
        1185 => x"13550701",
        1186 => x"b357f300",
        1187 => x"3318b300",
        1188 => x"33d3a602",
        1189 => x"13160701",
        1190 => x"b398b800",
        1191 => x"13560601",
        1192 => x"b3e71701",
        1193 => x"b3f6a602",
        1194 => x"b3086602",
        1195 => x"93950601",
        1196 => x"93d60701",
        1197 => x"b3e6b600",
        1198 => x"93050300",
        1199 => x"63fe1601",
        1200 => x"b386e600",
        1201 => x"9305f3ff",
        1202 => x"63e8e600",
        1203 => x"63f61601",
        1204 => x"9305e3ff",
        1205 => x"b386e600",
        1206 => x"b3861641",
        1207 => x"b3d8a602",
        1208 => x"93970701",
        1209 => x"93d70701",
        1210 => x"b3f6a602",
        1211 => x"33061603",
        1212 => x"93960601",
        1213 => x"b3e7d700",
        1214 => x"93860800",
        1215 => x"63fec700",
        1216 => x"b387e700",
        1217 => x"9386f8ff",
        1218 => x"63e8e700",
        1219 => x"63f6c700",
        1220 => x"9386e8ff",
        1221 => x"b387e700",
        1222 => x"93950501",
        1223 => x"b387c740",
        1224 => x"b3e5d500",
        1225 => x"6ff09feb",
        1226 => x"63e6d518",
        1227 => x"b7070100",
        1228 => x"63f4f604",
        1229 => x"13b70610",
        1230 => x"13471700",
        1231 => x"13173700",
        1232 => x"b7370000",
        1233 => x"b3d5e600",
        1234 => x"9387470e",
        1235 => x"b387b700",
        1236 => x"83c70700",
        1237 => x"b387e700",
        1238 => x"13070002",
        1239 => x"b305f740",
        1240 => x"6316f702",
        1241 => x"13051000",
        1242 => x"e3ee16e1",
        1243 => x"3335c300",
        1244 => x"13451500",
        1245 => x"67800000",
        1246 => x"b7070001",
        1247 => x"13070001",
        1248 => x"e3e0f6fc",
        1249 => x"13078001",
        1250 => x"6ff09ffb",
        1251 => x"3357f600",
        1252 => x"b396b600",
        1253 => x"b366d700",
        1254 => x"33d7f800",
        1255 => x"b398b800",
        1256 => x"b357f300",
        1257 => x"b3e71701",
        1258 => x"93d80601",
        1259 => x"b35e1703",
        1260 => x"13980601",
        1261 => x"13580801",
        1262 => x"3316b600",
        1263 => x"33771703",
        1264 => x"330ed803",
        1265 => x"13150701",
        1266 => x"13d70701",
        1267 => x"3367a700",
        1268 => x"13850e00",
        1269 => x"637ec701",
        1270 => x"3307d700",
        1271 => x"1385feff",
        1272 => x"6368d700",
        1273 => x"6376c701",
        1274 => x"1385eeff",
        1275 => x"3307d700",
        1276 => x"3307c741",
        1277 => x"335e1703",
        1278 => x"93970701",
        1279 => x"93d70701",
        1280 => x"33771703",
        1281 => x"3308c803",
        1282 => x"13170701",
        1283 => x"b3e7e700",
        1284 => x"13070e00",
        1285 => x"63fe0701",
        1286 => x"b387d700",
        1287 => x"1307feff",
        1288 => x"63e8d700",
        1289 => x"63f60701",
        1290 => x"1307eeff",
        1291 => x"b387d700",
        1292 => x"13150501",
        1293 => x"370e0100",
        1294 => x"3365e500",
        1295 => x"9306feff",
        1296 => x"3377d500",
        1297 => x"b3870741",
        1298 => x"b376d600",
        1299 => x"13580501",
        1300 => x"13560601",
        1301 => x"b308d702",
        1302 => x"b306d802",
        1303 => x"3307c702",
        1304 => x"3308c802",
        1305 => x"3306d700",
        1306 => x"13d70801",
        1307 => x"3307c700",
        1308 => x"6374d700",
        1309 => x"3308c801",
        1310 => x"93560701",
        1311 => x"b3860601",
        1312 => x"63e6d702",
        1313 => x"e39ed7ce",
        1314 => x"b7070100",
        1315 => x"9387f7ff",
        1316 => x"3377f700",
        1317 => x"13170701",
        1318 => x"b3f8f800",
        1319 => x"3313b300",
        1320 => x"33071701",
        1321 => x"93050000",
        1322 => x"e37ee3cc",
        1323 => x"1305f5ff",
        1324 => x"6ff01fcd",
        1325 => x"93050000",
        1326 => x"13050000",
        1327 => x"67800000",
        1328 => x"13080600",
        1329 => x"93070500",
        1330 => x"13870500",
        1331 => x"63960620",
        1332 => x"b7380000",
        1333 => x"9388480e",
        1334 => x"63fcc50c",
        1335 => x"b7060100",
        1336 => x"637ed60a",
        1337 => x"93360610",
        1338 => x"93c61600",
        1339 => x"93963600",
        1340 => x"3353d600",
        1341 => x"b3886800",
        1342 => x"83c80800",
        1343 => x"13030002",
        1344 => x"b386d800",
        1345 => x"b308d340",
        1346 => x"630cd300",
        1347 => x"33971501",
        1348 => x"b356d500",
        1349 => x"33181601",
        1350 => x"33e7e600",
        1351 => x"b3171501",
        1352 => x"13560801",
        1353 => x"b356c702",
        1354 => x"13150801",
        1355 => x"13550501",
        1356 => x"3377c702",
        1357 => x"b386a602",
        1358 => x"93150701",
        1359 => x"13d70701",
        1360 => x"3367b700",
        1361 => x"637ad700",
        1362 => x"33070701",
        1363 => x"63660701",
        1364 => x"6374d700",
        1365 => x"33070701",
        1366 => x"3307d740",
        1367 => x"b356c702",
        1368 => x"3377c702",
        1369 => x"b386a602",
        1370 => x"93970701",
        1371 => x"13170701",
        1372 => x"93d70701",
        1373 => x"b3e7e700",
        1374 => x"63fad700",
        1375 => x"b3870701",
        1376 => x"63e60701",
        1377 => x"63f4d700",
        1378 => x"b3870701",
        1379 => x"b387d740",
        1380 => x"33d51701",
        1381 => x"93050000",
        1382 => x"67800000",
        1383 => x"37030001",
        1384 => x"93060001",
        1385 => x"e36666f4",
        1386 => x"93068001",
        1387 => x"6ff05ff4",
        1388 => x"63140600",
        1389 => x"73001000",
        1390 => x"37070100",
        1391 => x"637ee606",
        1392 => x"93360610",
        1393 => x"93c61600",
        1394 => x"93963600",
        1395 => x"3357d600",
        1396 => x"b388e800",
        1397 => x"03c70800",
        1398 => x"3307d700",
        1399 => x"93060002",
        1400 => x"b388e640",
        1401 => x"6394e606",
        1402 => x"3387c540",
        1403 => x"93550801",
        1404 => x"3356b702",
        1405 => x"13150801",
        1406 => x"13550501",
        1407 => x"93d60701",
        1408 => x"3377b702",
        1409 => x"3306a602",
        1410 => x"13170701",
        1411 => x"33e7e600",
        1412 => x"637ac700",
        1413 => x"33070701",
        1414 => x"63660701",
        1415 => x"6374c700",
        1416 => x"33070701",
        1417 => x"3307c740",
        1418 => x"b356b702",
        1419 => x"3377b702",
        1420 => x"b386a602",
        1421 => x"6ff05ff3",
        1422 => x"37070001",
        1423 => x"93060001",
        1424 => x"e366e6f8",
        1425 => x"93068001",
        1426 => x"6ff05ff8",
        1427 => x"33181601",
        1428 => x"b3d6e500",
        1429 => x"b3171501",
        1430 => x"b3951501",
        1431 => x"3357e500",
        1432 => x"13550801",
        1433 => x"3367b700",
        1434 => x"b3d5a602",
        1435 => x"13130801",
        1436 => x"13530301",
        1437 => x"b3f6a602",
        1438 => x"b3856502",
        1439 => x"13960601",
        1440 => x"93560701",
        1441 => x"b3e6c600",
        1442 => x"63fab600",
        1443 => x"b3860601",
        1444 => x"63e60601",
        1445 => x"63f4b600",
        1446 => x"b3860601",
        1447 => x"b386b640",
        1448 => x"33d6a602",
        1449 => x"13170701",
        1450 => x"13570701",
        1451 => x"b3f6a602",
        1452 => x"33066602",
        1453 => x"93960601",
        1454 => x"3367d700",
        1455 => x"637ac700",
        1456 => x"33070701",
        1457 => x"63660701",
        1458 => x"6374c700",
        1459 => x"33070701",
        1460 => x"3307c740",
        1461 => x"6ff09ff1",
        1462 => x"63e4d51c",
        1463 => x"37080100",
        1464 => x"63fe0605",
        1465 => x"13b80610",
        1466 => x"13481800",
        1467 => x"13183800",
        1468 => x"b7380000",
        1469 => x"33d30601",
        1470 => x"9388480e",
        1471 => x"b3886800",
        1472 => x"83c80800",
        1473 => x"13030002",
        1474 => x"b3880801",
        1475 => x"33081341",
        1476 => x"63101305",
        1477 => x"63e4b600",
        1478 => x"636cc500",
        1479 => x"3306c540",
        1480 => x"b386d540",
        1481 => x"3337c500",
        1482 => x"3387e640",
        1483 => x"93070600",
        1484 => x"13850700",
        1485 => x"93050700",
        1486 => x"67800000",
        1487 => x"b7080001",
        1488 => x"13080001",
        1489 => x"e3e616fb",
        1490 => x"13088001",
        1491 => x"6ff05ffa",
        1492 => x"b3960601",
        1493 => x"33531601",
        1494 => x"3363d300",
        1495 => x"135e0301",
        1496 => x"b3d61501",
        1497 => x"33dfc603",
        1498 => x"13170301",
        1499 => x"13570701",
        1500 => x"b3970501",
        1501 => x"b3551501",
        1502 => x"b3e5f500",
        1503 => x"93d70501",
        1504 => x"33160601",
        1505 => x"33150501",
        1506 => x"b3f6c603",
        1507 => x"b30ee703",
        1508 => x"93960601",
        1509 => x"b3e7d700",
        1510 => x"93060f00",
        1511 => x"63fed701",
        1512 => x"b3876700",
        1513 => x"9306ffff",
        1514 => x"63e86700",
        1515 => x"63f6d701",
        1516 => x"9306efff",
        1517 => x"b3876700",
        1518 => x"b387d741",
        1519 => x"b3dec703",
        1520 => x"93950501",
        1521 => x"93d50501",
        1522 => x"b3f7c703",
        1523 => x"3307d703",
        1524 => x"93970701",
        1525 => x"b3e5f500",
        1526 => x"93870e00",
        1527 => x"63fee500",
        1528 => x"b3856500",
        1529 => x"9387feff",
        1530 => x"63e86500",
        1531 => x"63f6e500",
        1532 => x"9387eeff",
        1533 => x"b3856500",
        1534 => x"93960601",
        1535 => x"370f0100",
        1536 => x"b3e6f600",
        1537 => x"9307ffff",
        1538 => x"135e0601",
        1539 => x"b385e540",
        1540 => x"33f7f600",
        1541 => x"93d60601",
        1542 => x"b377f600",
        1543 => x"b30ef702",
        1544 => x"b387f602",
        1545 => x"3307c703",
        1546 => x"b386c603",
        1547 => x"330ef700",
        1548 => x"13d70e01",
        1549 => x"3307c701",
        1550 => x"6374f700",
        1551 => x"b386e601",
        1552 => x"93570701",
        1553 => x"b387d700",
        1554 => x"b7060100",
        1555 => x"9386f6ff",
        1556 => x"3377d700",
        1557 => x"13170701",
        1558 => x"b3fede00",
        1559 => x"3307d701",
        1560 => x"63e6f500",
        1561 => x"639ef500",
        1562 => x"637ce500",
        1563 => x"3306c740",
        1564 => x"3337c700",
        1565 => x"33076700",
        1566 => x"b387e740",
        1567 => x"13070600",
        1568 => x"3307e540",
        1569 => x"3335e500",
        1570 => x"b385f540",
        1571 => x"b385a540",
        1572 => x"b3981501",
        1573 => x"33570701",
        1574 => x"33e5e800",
        1575 => x"b3d50501",
        1576 => x"67800000",
        1577 => x"13030500",
        1578 => x"630e0600",
        1579 => x"83830500",
        1580 => x"23007300",
        1581 => x"1306f6ff",
        1582 => x"13031300",
        1583 => x"93851500",
        1584 => x"e31606fe",
        1585 => x"67800000",
        1586 => x"13030500",
        1587 => x"630a0600",
        1588 => x"2300b300",
        1589 => x"1306f6ff",
        1590 => x"13031300",
        1591 => x"e31a06fe",
        1592 => x"67800000",
        1593 => x"630c0602",
        1594 => x"13030500",
        1595 => x"93061000",
        1596 => x"636ab500",
        1597 => x"9306f0ff",
        1598 => x"1307f6ff",
        1599 => x"3303e300",
        1600 => x"b385e500",
        1601 => x"83830500",
        1602 => x"23007300",
        1603 => x"1306f6ff",
        1604 => x"3303d300",
        1605 => x"b385d500",
        1606 => x"e31606fe",
        1607 => x"67800000",
        1608 => x"130101f9",
        1609 => x"23248106",
        1610 => x"232e3105",
        1611 => x"23261106",
        1612 => x"23229106",
        1613 => x"23202107",
        1614 => x"232c4105",
        1615 => x"232a5105",
        1616 => x"23286105",
        1617 => x"23267105",
        1618 => x"23248105",
        1619 => x"93090500",
        1620 => x"13840500",
        1621 => x"232c0100",
        1622 => x"232e0100",
        1623 => x"23200102",
        1624 => x"23220102",
        1625 => x"23240102",
        1626 => x"23260102",
        1627 => x"23280102",
        1628 => x"232a0102",
        1629 => x"232c0102",
        1630 => x"232e0102",
        1631 => x"97f2ffff",
        1632 => x"93828295",
        1633 => x"73905230",
        1634 => x"73e05030",
        1635 => x"b7220000",
        1636 => x"93828280",
        1637 => x"73900230",
        1638 => x"efe04fee",
        1639 => x"b7877d01",
        1640 => x"370700f0",
        1641 => x"9387f783",
        1642 => x"2326f708",
        1643 => x"37390000",
        1644 => x"93071001",
        1645 => x"2320f708",
        1646 => x"13050921",
        1647 => x"efe0cfef",
        1648 => x"63543003",
        1649 => x"9384f9ff",
        1650 => x"9309f0ff",
        1651 => x"03250400",
        1652 => x"9384f4ff",
        1653 => x"13044400",
        1654 => x"efe00fee",
        1655 => x"13050921",
        1656 => x"efe08fed",
        1657 => x"e39434ff",
        1658 => x"37350000",
        1659 => x"1305451e",
        1660 => x"371a0000",
        1661 => x"efe04fec",
        1662 => x"13040000",
        1663 => x"373c0000",
        1664 => x"130a0ae1",
        1665 => x"930a0000",
        1666 => x"930b0019",
        1667 => x"93050000",
        1668 => x"13058100",
        1669 => x"ef00c026",
        1670 => x"13041400",
        1671 => x"63020502",
        1672 => x"e31674ff",
        1673 => x"73001000",
        1674 => x"93050000",
        1675 => x"13058100",
        1676 => x"13040000",
        1677 => x"ef00c024",
        1678 => x"13041400",
        1679 => x"e31205fe",
        1680 => x"83248100",
        1681 => x"032bc100",
        1682 => x"1306c003",
        1683 => x"93060000",
        1684 => x"13850400",
        1685 => x"93050b00",
        1686 => x"eff08f9e",
        1687 => x"93090500",
        1688 => x"1306c003",
        1689 => x"93060000",
        1690 => x"13850400",
        1691 => x"93050b00",
        1692 => x"efe09fd5",
        1693 => x"1306c003",
        1694 => x"93060000",
        1695 => x"eff04f9c",
        1696 => x"13060a00",
        1697 => x"93860a00",
        1698 => x"13090500",
        1699 => x"93050b00",
        1700 => x"13850400",
        1701 => x"efe05fd3",
        1702 => x"83260101",
        1703 => x"13070500",
        1704 => x"13880900",
        1705 => x"93070900",
        1706 => x"13860400",
        1707 => x"93054c21",
        1708 => x"13058101",
        1709 => x"ef00c015",
        1710 => x"13058101",
        1711 => x"efe0cfdf",
        1712 => x"e31674f5",
        1713 => x"6ff01ff6",
        1714 => x"03a5c187",
        1715 => x"67800000",
        1716 => x"130101ff",
        1717 => x"23248100",
        1718 => x"23261100",
        1719 => x"93070000",
        1720 => x"13040500",
        1721 => x"63880700",
        1722 => x"93050000",
        1723 => x"97000000",
        1724 => x"e7000000",
        1725 => x"b7370000",
        1726 => x"03a54738",
        1727 => x"83278502",
        1728 => x"63840700",
        1729 => x"e7800700",
        1730 => x"13050400",
        1731 => x"ef108033",
        1732 => x"130101ff",
        1733 => x"23248100",
        1734 => x"23229100",
        1735 => x"37340000",
        1736 => x"b7340000",
        1737 => x"93878438",
        1738 => x"13048438",
        1739 => x"3304f440",
        1740 => x"23202101",
        1741 => x"23261100",
        1742 => x"13542440",
        1743 => x"93848438",
        1744 => x"13090000",
        1745 => x"63108904",
        1746 => x"b7340000",
        1747 => x"37340000",
        1748 => x"93878438",
        1749 => x"13048438",
        1750 => x"3304f440",
        1751 => x"13542440",
        1752 => x"93848438",
        1753 => x"13090000",
        1754 => x"63188902",
        1755 => x"8320c100",
        1756 => x"03248100",
        1757 => x"83244100",
        1758 => x"03290100",
        1759 => x"13010101",
        1760 => x"67800000",
        1761 => x"83a70400",
        1762 => x"13091900",
        1763 => x"93844400",
        1764 => x"e7800700",
        1765 => x"6ff01ffb",
        1766 => x"83a70400",
        1767 => x"13091900",
        1768 => x"93844400",
        1769 => x"e7800700",
        1770 => x"6ff01ffc",
        1771 => x"130101f6",
        1772 => x"232af108",
        1773 => x"b7070080",
        1774 => x"93c7f7ff",
        1775 => x"232ef100",
        1776 => x"2328f100",
        1777 => x"b707ffff",
        1778 => x"2326d108",
        1779 => x"2324b100",
        1780 => x"232cb100",
        1781 => x"93878720",
        1782 => x"9306c108",
        1783 => x"93058100",
        1784 => x"232e1106",
        1785 => x"232af100",
        1786 => x"2328e108",
        1787 => x"232c0109",
        1788 => x"232e1109",
        1789 => x"2322d100",
        1790 => x"ef004041",
        1791 => x"83278100",
        1792 => x"23800700",
        1793 => x"8320c107",
        1794 => x"1301010a",
        1795 => x"67800000",
        1796 => x"130101f6",
        1797 => x"232af108",
        1798 => x"b7070080",
        1799 => x"93c7f7ff",
        1800 => x"232ef100",
        1801 => x"2328f100",
        1802 => x"b707ffff",
        1803 => x"93878720",
        1804 => x"232af100",
        1805 => x"2324a100",
        1806 => x"232ca100",
        1807 => x"03a5c187",
        1808 => x"2324c108",
        1809 => x"2326d108",
        1810 => x"13860500",
        1811 => x"93068108",
        1812 => x"93058100",
        1813 => x"232e1106",
        1814 => x"2328e108",
        1815 => x"232c0109",
        1816 => x"232e1109",
        1817 => x"2322d100",
        1818 => x"ef00403a",
        1819 => x"83278100",
        1820 => x"23800700",
        1821 => x"8320c107",
        1822 => x"1301010a",
        1823 => x"67800000",
        1824 => x"13860500",
        1825 => x"93050500",
        1826 => x"03a5c187",
        1827 => x"6f004000",
        1828 => x"130101ff",
        1829 => x"23248100",
        1830 => x"23229100",
        1831 => x"13040500",
        1832 => x"13850500",
        1833 => x"93050600",
        1834 => x"23261100",
        1835 => x"23a20188",
        1836 => x"ef10401c",
        1837 => x"9307f0ff",
        1838 => x"6318f500",
        1839 => x"83a74188",
        1840 => x"63840700",
        1841 => x"2320f400",
        1842 => x"8320c100",
        1843 => x"03248100",
        1844 => x"83244100",
        1845 => x"13010101",
        1846 => x"67800000",
        1847 => x"130101fe",
        1848 => x"23282101",
        1849 => x"03a98500",
        1850 => x"232c8100",
        1851 => x"23263101",
        1852 => x"23244101",
        1853 => x"23225101",
        1854 => x"232e1100",
        1855 => x"232a9100",
        1856 => x"23206101",
        1857 => x"83aa0500",
        1858 => x"13840500",
        1859 => x"130a0600",
        1860 => x"93890600",
        1861 => x"63ec2609",
        1862 => x"83d7c500",
        1863 => x"13f70748",
        1864 => x"63040708",
        1865 => x"03274401",
        1866 => x"93043000",
        1867 => x"83a50501",
        1868 => x"b384e402",
        1869 => x"13072000",
        1870 => x"b38aba40",
        1871 => x"130b0500",
        1872 => x"b3c4e402",
        1873 => x"13871600",
        1874 => x"33075701",
        1875 => x"63f4e400",
        1876 => x"93040700",
        1877 => x"93f70740",
        1878 => x"6386070a",
        1879 => x"93850400",
        1880 => x"13050b00",
        1881 => x"ef001065",
        1882 => x"13090500",
        1883 => x"630c050a",
        1884 => x"83250401",
        1885 => x"13860a00",
        1886 => x"eff0dfb2",
        1887 => x"8357c400",
        1888 => x"93f7f7b7",
        1889 => x"93e70708",
        1890 => x"2316f400",
        1891 => x"23282401",
        1892 => x"232a9400",
        1893 => x"33095901",
        1894 => x"b3845441",
        1895 => x"23202401",
        1896 => x"23249400",
        1897 => x"13890900",
        1898 => x"63f42901",
        1899 => x"13890900",
        1900 => x"03250400",
        1901 => x"13060900",
        1902 => x"93050a00",
        1903 => x"eff09fb2",
        1904 => x"83278400",
        1905 => x"13050000",
        1906 => x"b3872741",
        1907 => x"2324f400",
        1908 => x"83270400",
        1909 => x"b3872701",
        1910 => x"2320f400",
        1911 => x"8320c101",
        1912 => x"03248101",
        1913 => x"83244101",
        1914 => x"03290101",
        1915 => x"8329c100",
        1916 => x"032a8100",
        1917 => x"832a4100",
        1918 => x"032b0100",
        1919 => x"13010102",
        1920 => x"67800000",
        1921 => x"13860400",
        1922 => x"13050b00",
        1923 => x"ef00906f",
        1924 => x"13090500",
        1925 => x"e31c05f6",
        1926 => x"83250401",
        1927 => x"13050b00",
        1928 => x"ef00d049",
        1929 => x"9307c000",
        1930 => x"2320fb00",
        1931 => x"8357c400",
        1932 => x"1305f0ff",
        1933 => x"93e70704",
        1934 => x"2316f400",
        1935 => x"6ff01ffa",
        1936 => x"83278600",
        1937 => x"130101fd",
        1938 => x"232e3101",
        1939 => x"23286101",
        1940 => x"23261102",
        1941 => x"23248102",
        1942 => x"23229102",
        1943 => x"23202103",
        1944 => x"232c4101",
        1945 => x"232a5101",
        1946 => x"23267101",
        1947 => x"23248101",
        1948 => x"23229101",
        1949 => x"2320a101",
        1950 => x"032b0600",
        1951 => x"93090600",
        1952 => x"63980712",
        1953 => x"13050000",
        1954 => x"8320c102",
        1955 => x"03248102",
        1956 => x"23a20900",
        1957 => x"83244102",
        1958 => x"03290102",
        1959 => x"8329c101",
        1960 => x"032a8101",
        1961 => x"832a4101",
        1962 => x"032b0101",
        1963 => x"832bc100",
        1964 => x"032c8100",
        1965 => x"832c4100",
        1966 => x"032d0100",
        1967 => x"13010103",
        1968 => x"67800000",
        1969 => x"832a0b00",
        1970 => x"032d4b00",
        1971 => x"130b8b00",
        1972 => x"03298400",
        1973 => x"832c0400",
        1974 => x"e3060dfe",
        1975 => x"63642d09",
        1976 => x"8357c400",
        1977 => x"13f70748",
        1978 => x"630e0706",
        1979 => x"83244401",
        1980 => x"83250401",
        1981 => x"b3849b02",
        1982 => x"b38cbc40",
        1983 => x"13871c00",
        1984 => x"3307a701",
        1985 => x"b3c48403",
        1986 => x"63f4e400",
        1987 => x"93040700",
        1988 => x"93f70740",
        1989 => x"638c070a",
        1990 => x"93850400",
        1991 => x"13050a00",
        1992 => x"ef005049",
        1993 => x"13090500",
        1994 => x"6302050c",
        1995 => x"83250401",
        1996 => x"13860c00",
        1997 => x"eff01f97",
        1998 => x"8357c400",
        1999 => x"93f7f7b7",
        2000 => x"93e70708",
        2001 => x"2316f400",
        2002 => x"23282401",
        2003 => x"232a9400",
        2004 => x"33099901",
        2005 => x"b3849441",
        2006 => x"23202401",
        2007 => x"23249400",
        2008 => x"13090d00",
        2009 => x"63742d01",
        2010 => x"13090d00",
        2011 => x"03250400",
        2012 => x"93850a00",
        2013 => x"13060900",
        2014 => x"eff0df96",
        2015 => x"83278400",
        2016 => x"b38aaa01",
        2017 => x"b3872741",
        2018 => x"2324f400",
        2019 => x"83270400",
        2020 => x"b3872701",
        2021 => x"2320f400",
        2022 => x"83a78900",
        2023 => x"b387a741",
        2024 => x"23a4f900",
        2025 => x"e38007ee",
        2026 => x"130d0000",
        2027 => x"6ff05ff2",
        2028 => x"130a0500",
        2029 => x"13840500",
        2030 => x"930a0000",
        2031 => x"130d0000",
        2032 => x"930b3000",
        2033 => x"130c2000",
        2034 => x"6ff09ff0",
        2035 => x"13860400",
        2036 => x"13050a00",
        2037 => x"ef001053",
        2038 => x"13090500",
        2039 => x"e31605f6",
        2040 => x"83250401",
        2041 => x"13050a00",
        2042 => x"ef00502d",
        2043 => x"9307c000",
        2044 => x"2320fa00",
        2045 => x"8357c400",
        2046 => x"1305f0ff",
        2047 => x"93e70704",
        2048 => x"2316f400",
        2049 => x"23a40900",
        2050 => x"6ff01fe8",
        2051 => x"83d7c500",
        2052 => x"130101f5",
        2053 => x"2324810a",
        2054 => x"2322910a",
        2055 => x"2320210b",
        2056 => x"232c4109",
        2057 => x"2326110a",
        2058 => x"232e3109",
        2059 => x"232a5109",
        2060 => x"23286109",
        2061 => x"23267109",
        2062 => x"23248109",
        2063 => x"23229109",
        2064 => x"2320a109",
        2065 => x"232eb107",
        2066 => x"93f70708",
        2067 => x"130a0500",
        2068 => x"13890500",
        2069 => x"93040600",
        2070 => x"13840600",
        2071 => x"63880706",
        2072 => x"83a70501",
        2073 => x"63940706",
        2074 => x"93050004",
        2075 => x"ef009034",
        2076 => x"2320a900",
        2077 => x"2328a900",
        2078 => x"63160504",
        2079 => x"9307c000",
        2080 => x"2320fa00",
        2081 => x"1305f0ff",
        2082 => x"8320c10a",
        2083 => x"0324810a",
        2084 => x"8324410a",
        2085 => x"0329010a",
        2086 => x"8329c109",
        2087 => x"032a8109",
        2088 => x"832a4109",
        2089 => x"032b0109",
        2090 => x"832bc108",
        2091 => x"032c8108",
        2092 => x"832c4108",
        2093 => x"032d0108",
        2094 => x"832dc107",
        2095 => x"1301010b",
        2096 => x"67800000",
        2097 => x"93070004",
        2098 => x"232af900",
        2099 => x"93070002",
        2100 => x"a304f102",
        2101 => x"93070003",
        2102 => x"23220102",
        2103 => x"2305f102",
        2104 => x"23268100",
        2105 => x"930c5002",
        2106 => x"373b0000",
        2107 => x"b73b0000",
        2108 => x"373d0000",
        2109 => x"372c0000",
        2110 => x"930a0000",
        2111 => x"13840400",
        2112 => x"83470400",
        2113 => x"63840700",
        2114 => x"639c970d",
        2115 => x"b30d9440",
        2116 => x"63069402",
        2117 => x"93860d00",
        2118 => x"13860400",
        2119 => x"93050900",
        2120 => x"13050a00",
        2121 => x"eff09fbb",
        2122 => x"9307f0ff",
        2123 => x"6306f524",
        2124 => x"83274102",
        2125 => x"b387b701",
        2126 => x"2322f102",
        2127 => x"83470400",
        2128 => x"638c0722",
        2129 => x"9307f0ff",
        2130 => x"93041400",
        2131 => x"23280100",
        2132 => x"232e0100",
        2133 => x"232af100",
        2134 => x"232c0100",
        2135 => x"a3090104",
        2136 => x"23240106",
        2137 => x"930d1000",
        2138 => x"83c50400",
        2139 => x"13065000",
        2140 => x"13050b2f",
        2141 => x"ef005012",
        2142 => x"83270101",
        2143 => x"13841400",
        2144 => x"63140506",
        2145 => x"13f70701",
        2146 => x"63060700",
        2147 => x"13070002",
        2148 => x"a309e104",
        2149 => x"13f78700",
        2150 => x"63060700",
        2151 => x"1307b002",
        2152 => x"a309e104",
        2153 => x"83c60400",
        2154 => x"1307a002",
        2155 => x"638ce604",
        2156 => x"8327c101",
        2157 => x"13840400",
        2158 => x"93060000",
        2159 => x"13069000",
        2160 => x"1305a000",
        2161 => x"03470400",
        2162 => x"93051400",
        2163 => x"130707fd",
        2164 => x"637ce608",
        2165 => x"63840604",
        2166 => x"232ef100",
        2167 => x"6f000004",
        2168 => x"13041400",
        2169 => x"6ff0dff1",
        2170 => x"13070b2f",
        2171 => x"3305e540",
        2172 => x"3395ad00",
        2173 => x"b3e7a700",
        2174 => x"2328f100",
        2175 => x"93040400",
        2176 => x"6ff09ff6",
        2177 => x"0327c100",
        2178 => x"93064700",
        2179 => x"03270700",
        2180 => x"2326d100",
        2181 => x"63400704",
        2182 => x"232ee100",
        2183 => x"03470400",
        2184 => x"9307e002",
        2185 => x"6316f708",
        2186 => x"03471400",
        2187 => x"9307a002",
        2188 => x"631af704",
        2189 => x"8327c100",
        2190 => x"13042400",
        2191 => x"13874700",
        2192 => x"83a70700",
        2193 => x"2326e100",
        2194 => x"63ca0702",
        2195 => x"232af100",
        2196 => x"6f000006",
        2197 => x"3307e040",
        2198 => x"93e72700",
        2199 => x"232ee100",
        2200 => x"2328f100",
        2201 => x"6ff09ffb",
        2202 => x"b387a702",
        2203 => x"13840500",
        2204 => x"93061000",
        2205 => x"b387e700",
        2206 => x"6ff0dff4",
        2207 => x"9307f0ff",
        2208 => x"6ff0dffc",
        2209 => x"13041400",
        2210 => x"232a0100",
        2211 => x"93060000",
        2212 => x"93070000",
        2213 => x"13069000",
        2214 => x"1305a000",
        2215 => x"03470400",
        2216 => x"93051400",
        2217 => x"130707fd",
        2218 => x"6372e608",
        2219 => x"e39006fa",
        2220 => x"83450400",
        2221 => x"13063000",
        2222 => x"13858b2f",
        2223 => x"ef00c07d",
        2224 => x"63020502",
        2225 => x"93878b2f",
        2226 => x"3305f540",
        2227 => x"83270101",
        2228 => x"13070004",
        2229 => x"3317a700",
        2230 => x"b3e7e700",
        2231 => x"13041400",
        2232 => x"2328f100",
        2233 => x"83450400",
        2234 => x"13066000",
        2235 => x"1305cd2f",
        2236 => x"93041400",
        2237 => x"2304b102",
        2238 => x"ef00007a",
        2239 => x"630a0508",
        2240 => x"63980a04",
        2241 => x"03270101",
        2242 => x"8327c100",
        2243 => x"13770710",
        2244 => x"63080702",
        2245 => x"93874700",
        2246 => x"2326f100",
        2247 => x"83274102",
        2248 => x"b3873701",
        2249 => x"2322f102",
        2250 => x"6ff05fdd",
        2251 => x"b387a702",
        2252 => x"13840500",
        2253 => x"93061000",
        2254 => x"b387e700",
        2255 => x"6ff01ff6",
        2256 => x"93877700",
        2257 => x"93f787ff",
        2258 => x"93878700",
        2259 => x"6ff0dffc",
        2260 => x"1307c100",
        2261 => x"9306cccd",
        2262 => x"13060900",
        2263 => x"93050101",
        2264 => x"13050a00",
        2265 => x"97000000",
        2266 => x"e7000000",
        2267 => x"9307f0ff",
        2268 => x"93090500",
        2269 => x"e314f5fa",
        2270 => x"8357c900",
        2271 => x"1305f0ff",
        2272 => x"93f70704",
        2273 => x"e39207d0",
        2274 => x"03254102",
        2275 => x"6ff0dfcf",
        2276 => x"1307c100",
        2277 => x"9306cccd",
        2278 => x"13060900",
        2279 => x"93050101",
        2280 => x"13050a00",
        2281 => x"ef00801b",
        2282 => x"6ff05ffc",
        2283 => x"130101fd",
        2284 => x"232c4101",
        2285 => x"83a70501",
        2286 => x"130a0700",
        2287 => x"03a78500",
        2288 => x"23248102",
        2289 => x"23202103",
        2290 => x"232e3101",
        2291 => x"232a5101",
        2292 => x"23261102",
        2293 => x"23229102",
        2294 => x"23286101",
        2295 => x"23267101",
        2296 => x"93090500",
        2297 => x"13840500",
        2298 => x"13090600",
        2299 => x"938a0600",
        2300 => x"63d4e700",
        2301 => x"93070700",
        2302 => x"2320f900",
        2303 => x"03473404",
        2304 => x"63060700",
        2305 => x"93871700",
        2306 => x"2320f900",
        2307 => x"83270400",
        2308 => x"93f70702",
        2309 => x"63880700",
        2310 => x"83270900",
        2311 => x"93872700",
        2312 => x"2320f900",
        2313 => x"83240400",
        2314 => x"93f46400",
        2315 => x"639e0400",
        2316 => x"130b9401",
        2317 => x"930bf0ff",
        2318 => x"8327c400",
        2319 => x"03270900",
        2320 => x"b387e740",
        2321 => x"63c2f408",
        2322 => x"83473404",
        2323 => x"b336f000",
        2324 => x"83270400",
        2325 => x"93f70702",
        2326 => x"6390070c",
        2327 => x"13063404",
        2328 => x"93850a00",
        2329 => x"13850900",
        2330 => x"e7000a00",
        2331 => x"9307f0ff",
        2332 => x"6308f506",
        2333 => x"83270400",
        2334 => x"13074000",
        2335 => x"93040000",
        2336 => x"93f76700",
        2337 => x"639ce700",
        2338 => x"8324c400",
        2339 => x"83270900",
        2340 => x"b384f440",
        2341 => x"63d40400",
        2342 => x"93040000",
        2343 => x"83278400",
        2344 => x"03270401",
        2345 => x"6356f700",
        2346 => x"b387e740",
        2347 => x"b384f400",
        2348 => x"13090000",
        2349 => x"1304a401",
        2350 => x"130bf0ff",
        2351 => x"63902409",
        2352 => x"13050000",
        2353 => x"6f000002",
        2354 => x"93061000",
        2355 => x"13060b00",
        2356 => x"93850a00",
        2357 => x"13850900",
        2358 => x"e7000a00",
        2359 => x"631a7503",
        2360 => x"1305f0ff",
        2361 => x"8320c102",
        2362 => x"03248102",
        2363 => x"83244102",
        2364 => x"03290102",
        2365 => x"8329c101",
        2366 => x"032a8101",
        2367 => x"832a4101",
        2368 => x"032b0101",
        2369 => x"832bc100",
        2370 => x"13010103",
        2371 => x"67800000",
        2372 => x"93841400",
        2373 => x"6ff05ff2",
        2374 => x"3307d400",
        2375 => x"13060003",
        2376 => x"a301c704",
        2377 => x"03475404",
        2378 => x"93871600",
        2379 => x"b307f400",
        2380 => x"93862600",
        2381 => x"a381e704",
        2382 => x"6ff05ff2",
        2383 => x"93061000",
        2384 => x"13060400",
        2385 => x"93850a00",
        2386 => x"13850900",
        2387 => x"e7000a00",
        2388 => x"e30865f9",
        2389 => x"13091900",
        2390 => x"6ff05ff6",
        2391 => x"130101fd",
        2392 => x"23248102",
        2393 => x"23229102",
        2394 => x"23202103",
        2395 => x"232e3101",
        2396 => x"23261102",
        2397 => x"232c4101",
        2398 => x"232a5101",
        2399 => x"23286101",
        2400 => x"83c88501",
        2401 => x"93078007",
        2402 => x"93040500",
        2403 => x"13840500",
        2404 => x"13090600",
        2405 => x"93890600",
        2406 => x"63ee1701",
        2407 => x"93072006",
        2408 => x"93863504",
        2409 => x"63ee1701",
        2410 => x"63840828",
        2411 => x"93078005",
        2412 => x"6388f822",
        2413 => x"930a2404",
        2414 => x"23011405",
        2415 => x"6f004004",
        2416 => x"9387d8f9",
        2417 => x"93f7f70f",
        2418 => x"13065001",
        2419 => x"e364f6fe",
        2420 => x"37360000",
        2421 => x"93972700",
        2422 => x"1306c632",
        2423 => x"b387c700",
        2424 => x"83a70700",
        2425 => x"67800700",
        2426 => x"83270700",
        2427 => x"938a2504",
        2428 => x"93864700",
        2429 => x"83a70700",
        2430 => x"2320d700",
        2431 => x"2381f504",
        2432 => x"93071000",
        2433 => x"6f008026",
        2434 => x"83a70500",
        2435 => x"03250700",
        2436 => x"13f60708",
        2437 => x"93054500",
        2438 => x"63060602",
        2439 => x"83270500",
        2440 => x"2320b700",
        2441 => x"37380000",
        2442 => x"63d80700",
        2443 => x"1307d002",
        2444 => x"b307f040",
        2445 => x"a301e404",
        2446 => x"13084830",
        2447 => x"1307a000",
        2448 => x"6f008006",
        2449 => x"13f60704",
        2450 => x"83270500",
        2451 => x"2320b700",
        2452 => x"e30a06fc",
        2453 => x"93970701",
        2454 => x"93d70741",
        2455 => x"6ff09ffc",
        2456 => x"03a60500",
        2457 => x"83270700",
        2458 => x"13750608",
        2459 => x"93854700",
        2460 => x"63080500",
        2461 => x"2320b700",
        2462 => x"83a70700",
        2463 => x"6f004001",
        2464 => x"13760604",
        2465 => x"2320b700",
        2466 => x"e30806fe",
        2467 => x"83d70700",
        2468 => x"37380000",
        2469 => x"1307f006",
        2470 => x"13084830",
        2471 => x"6388e814",
        2472 => x"1307a000",
        2473 => x"a3010404",
        2474 => x"03264400",
        2475 => x"2324c400",
        2476 => x"63480600",
        2477 => x"83250400",
        2478 => x"93f5b5ff",
        2479 => x"2320b400",
        2480 => x"63960700",
        2481 => x"938a0600",
        2482 => x"63040602",
        2483 => x"938a0600",
        2484 => x"33f6e702",
        2485 => x"938afaff",
        2486 => x"3306c800",
        2487 => x"03460600",
        2488 => x"2380ca00",
        2489 => x"13860700",
        2490 => x"b3d7e702",
        2491 => x"e372e6fe",
        2492 => x"93078000",
        2493 => x"6314f702",
        2494 => x"83270400",
        2495 => x"93f71700",
        2496 => x"638e0700",
        2497 => x"03274400",
        2498 => x"83270401",
        2499 => x"63c8e700",
        2500 => x"93070003",
        2501 => x"a38ffafe",
        2502 => x"938afaff",
        2503 => x"b3865641",
        2504 => x"2328d400",
        2505 => x"13870900",
        2506 => x"93060900",
        2507 => x"1306c100",
        2508 => x"93050400",
        2509 => x"13850400",
        2510 => x"eff05fc7",
        2511 => x"130af0ff",
        2512 => x"631c4513",
        2513 => x"1305f0ff",
        2514 => x"8320c102",
        2515 => x"03248102",
        2516 => x"83244102",
        2517 => x"03290102",
        2518 => x"8329c101",
        2519 => x"032a8101",
        2520 => x"832a4101",
        2521 => x"032b0101",
        2522 => x"13010103",
        2523 => x"67800000",
        2524 => x"83a70500",
        2525 => x"93e70702",
        2526 => x"23a0f500",
        2527 => x"37380000",
        2528 => x"93088007",
        2529 => x"13088831",
        2530 => x"a3021405",
        2531 => x"03260400",
        2532 => x"83250700",
        2533 => x"13750608",
        2534 => x"83a70500",
        2535 => x"93854500",
        2536 => x"631a0500",
        2537 => x"13750604",
        2538 => x"63060500",
        2539 => x"93970701",
        2540 => x"93d70701",
        2541 => x"2320b700",
        2542 => x"13771600",
        2543 => x"63060700",
        2544 => x"13660602",
        2545 => x"2320c400",
        2546 => x"13070001",
        2547 => x"e39c07ec",
        2548 => x"03260400",
        2549 => x"1376f6fd",
        2550 => x"2320c400",
        2551 => x"6ff09fec",
        2552 => x"37380000",
        2553 => x"13084830",
        2554 => x"6ff01ffa",
        2555 => x"13078000",
        2556 => x"6ff05feb",
        2557 => x"03a60500",
        2558 => x"83270700",
        2559 => x"83a54501",
        2560 => x"13780608",
        2561 => x"13854700",
        2562 => x"630a0800",
        2563 => x"2320a700",
        2564 => x"83a70700",
        2565 => x"23a0b700",
        2566 => x"6f008001",
        2567 => x"2320a700",
        2568 => x"13760604",
        2569 => x"83a70700",
        2570 => x"e30606fe",
        2571 => x"2390b700",
        2572 => x"23280400",
        2573 => x"938a0600",
        2574 => x"6ff0dfee",
        2575 => x"83270700",
        2576 => x"03a64500",
        2577 => x"93050000",
        2578 => x"93864700",
        2579 => x"2320d700",
        2580 => x"83aa0700",
        2581 => x"13850a00",
        2582 => x"ef000024",
        2583 => x"63060500",
        2584 => x"33055541",
        2585 => x"2322a400",
        2586 => x"83274400",
        2587 => x"2328f400",
        2588 => x"a3010404",
        2589 => x"6ff01feb",
        2590 => x"83260401",
        2591 => x"13860a00",
        2592 => x"93050900",
        2593 => x"13850400",
        2594 => x"e7800900",
        2595 => x"e30c45eb",
        2596 => x"83270400",
        2597 => x"93f72700",
        2598 => x"63940704",
        2599 => x"8327c100",
        2600 => x"0325c400",
        2601 => x"e352f5ea",
        2602 => x"13850700",
        2603 => x"6ff0dfe9",
        2604 => x"93061000",
        2605 => x"13860a00",
        2606 => x"93050900",
        2607 => x"13850400",
        2608 => x"e7800900",
        2609 => x"e30065e9",
        2610 => x"130a1a00",
        2611 => x"8327c400",
        2612 => x"0327c100",
        2613 => x"b387e740",
        2614 => x"e34cfafc",
        2615 => x"6ff01ffc",
        2616 => x"130a0000",
        2617 => x"930a9401",
        2618 => x"130bf0ff",
        2619 => x"6ff01ffe",
        2620 => x"130101ff",
        2621 => x"23248100",
        2622 => x"13840500",
        2623 => x"83a50500",
        2624 => x"23229100",
        2625 => x"23261100",
        2626 => x"93040500",
        2627 => x"63840500",
        2628 => x"eff01ffe",
        2629 => x"93050400",
        2630 => x"03248100",
        2631 => x"8320c100",
        2632 => x"13850400",
        2633 => x"83244100",
        2634 => x"13010101",
        2635 => x"6f000019",
        2636 => x"83a7c187",
        2637 => x"6380a716",
        2638 => x"83274502",
        2639 => x"130101fe",
        2640 => x"232c8100",
        2641 => x"232e1100",
        2642 => x"232a9100",
        2643 => x"23282101",
        2644 => x"23263101",
        2645 => x"13040500",
        2646 => x"63840702",
        2647 => x"83a7c700",
        2648 => x"93040000",
        2649 => x"13090008",
        2650 => x"6392070e",
        2651 => x"83274402",
        2652 => x"83a50700",
        2653 => x"63860500",
        2654 => x"13050400",
        2655 => x"ef000014",
        2656 => x"83254401",
        2657 => x"63860500",
        2658 => x"13050400",
        2659 => x"ef000013",
        2660 => x"83254402",
        2661 => x"63860500",
        2662 => x"13050400",
        2663 => x"ef000012",
        2664 => x"83258403",
        2665 => x"63860500",
        2666 => x"13050400",
        2667 => x"ef000011",
        2668 => x"8325c403",
        2669 => x"63860500",
        2670 => x"13050400",
        2671 => x"ef000010",
        2672 => x"83250404",
        2673 => x"63860500",
        2674 => x"13050400",
        2675 => x"ef00000f",
        2676 => x"8325c405",
        2677 => x"63860500",
        2678 => x"13050400",
        2679 => x"ef00000e",
        2680 => x"83258405",
        2681 => x"63860500",
        2682 => x"13050400",
        2683 => x"ef00000d",
        2684 => x"83254403",
        2685 => x"63860500",
        2686 => x"13050400",
        2687 => x"ef00000c",
        2688 => x"83278401",
        2689 => x"638a0706",
        2690 => x"83278402",
        2691 => x"13050400",
        2692 => x"e7800700",
        2693 => x"83258404",
        2694 => x"63800506",
        2695 => x"13050400",
        2696 => x"03248101",
        2697 => x"8320c101",
        2698 => x"83244101",
        2699 => x"03290101",
        2700 => x"8329c100",
        2701 => x"13010102",
        2702 => x"6ff09feb",
        2703 => x"b3859500",
        2704 => x"83a50500",
        2705 => x"63900502",
        2706 => x"93844400",
        2707 => x"83274402",
        2708 => x"83a5c700",
        2709 => x"e39424ff",
        2710 => x"13050400",
        2711 => x"ef000006",
        2712 => x"6ff0dff0",
        2713 => x"83a90500",
        2714 => x"13050400",
        2715 => x"ef000005",
        2716 => x"93850900",
        2717 => x"6ff01ffd",
        2718 => x"8320c101",
        2719 => x"03248101",
        2720 => x"83244101",
        2721 => x"03290101",
        2722 => x"8329c100",
        2723 => x"13010102",
        2724 => x"67800000",
        2725 => x"67800000",
        2726 => x"93f5f50f",
        2727 => x"3306c500",
        2728 => x"6316c500",
        2729 => x"13050000",
        2730 => x"67800000",
        2731 => x"83470500",
        2732 => x"e38cb7fe",
        2733 => x"13051500",
        2734 => x"6ff09ffe",
        2735 => x"638a050e",
        2736 => x"83a7c5ff",
        2737 => x"130101fe",
        2738 => x"232c8100",
        2739 => x"232e1100",
        2740 => x"1384c5ff",
        2741 => x"63d40700",
        2742 => x"3304f400",
        2743 => x"2326a100",
        2744 => x"ef000034",
        2745 => x"83a78188",
        2746 => x"0325c100",
        2747 => x"639e0700",
        2748 => x"23220400",
        2749 => x"23a48188",
        2750 => x"03248101",
        2751 => x"8320c101",
        2752 => x"13010102",
        2753 => x"6f000032",
        2754 => x"6374f402",
        2755 => x"03260400",
        2756 => x"b306c400",
        2757 => x"639ad700",
        2758 => x"83a60700",
        2759 => x"83a74700",
        2760 => x"b386c600",
        2761 => x"2320d400",
        2762 => x"2322f400",
        2763 => x"6ff09ffc",
        2764 => x"13870700",
        2765 => x"83a74700",
        2766 => x"63840700",
        2767 => x"e37af4fe",
        2768 => x"83260700",
        2769 => x"3306d700",
        2770 => x"63188602",
        2771 => x"03260400",
        2772 => x"b386c600",
        2773 => x"2320d700",
        2774 => x"3306d700",
        2775 => x"e39ec7f8",
        2776 => x"03a60700",
        2777 => x"83a74700",
        2778 => x"b306d600",
        2779 => x"2320d700",
        2780 => x"2322f700",
        2781 => x"6ff05ff8",
        2782 => x"6378c400",
        2783 => x"9307c000",
        2784 => x"2320f500",
        2785 => x"6ff05ff7",
        2786 => x"03260400",
        2787 => x"b306c400",
        2788 => x"639ad700",
        2789 => x"83a60700",
        2790 => x"83a74700",
        2791 => x"b386c600",
        2792 => x"2320d400",
        2793 => x"2322f400",
        2794 => x"23228700",
        2795 => x"6ff0dff4",
        2796 => x"67800000",
        2797 => x"130101fe",
        2798 => x"232a9100",
        2799 => x"93843500",
        2800 => x"93f4c4ff",
        2801 => x"23282101",
        2802 => x"232e1100",
        2803 => x"232c8100",
        2804 => x"23263101",
        2805 => x"93848400",
        2806 => x"9307c000",
        2807 => x"13090500",
        2808 => x"63f4f406",
        2809 => x"9304c000",
        2810 => x"63e2b406",
        2811 => x"13050900",
        2812 => x"ef000023",
        2813 => x"03a78188",
        2814 => x"93868188",
        2815 => x"13040700",
        2816 => x"631a0406",
        2817 => x"1384c188",
        2818 => x"83270400",
        2819 => x"639a0700",
        2820 => x"93050000",
        2821 => x"13050900",
        2822 => x"ef00001c",
        2823 => x"2320a400",
        2824 => x"93850400",
        2825 => x"13050900",
        2826 => x"ef00001b",
        2827 => x"9309f0ff",
        2828 => x"631a350b",
        2829 => x"9307c000",
        2830 => x"2320f900",
        2831 => x"13050900",
        2832 => x"ef00401e",
        2833 => x"6f000001",
        2834 => x"e3d004fa",
        2835 => x"9307c000",
        2836 => x"2320f900",
        2837 => x"13050000",
        2838 => x"8320c101",
        2839 => x"03248101",
        2840 => x"83244101",
        2841 => x"03290101",
        2842 => x"8329c100",
        2843 => x"13010102",
        2844 => x"67800000",
        2845 => x"83270400",
        2846 => x"b3879740",
        2847 => x"63ce0704",
        2848 => x"1306b000",
        2849 => x"637af600",
        2850 => x"2320f400",
        2851 => x"3304f400",
        2852 => x"23209400",
        2853 => x"6f000001",
        2854 => x"83274400",
        2855 => x"631a8702",
        2856 => x"23a0f600",
        2857 => x"13050900",
        2858 => x"ef00c017",
        2859 => x"1305b400",
        2860 => x"93074400",
        2861 => x"137585ff",
        2862 => x"3307f540",
        2863 => x"e30ef5f8",
        2864 => x"3304e400",
        2865 => x"b387a740",
        2866 => x"2320f400",
        2867 => x"6ff0dff8",
        2868 => x"2322f700",
        2869 => x"6ff01ffd",
        2870 => x"13070400",
        2871 => x"03244400",
        2872 => x"6ff01ff2",
        2873 => x"13043500",
        2874 => x"1374c4ff",
        2875 => x"e30285fa",
        2876 => x"b305a440",
        2877 => x"13050900",
        2878 => x"ef00000e",
        2879 => x"e31a35f9",
        2880 => x"6ff05ff3",
        2881 => x"130101fe",
        2882 => x"232c8100",
        2883 => x"232e1100",
        2884 => x"232a9100",
        2885 => x"23282101",
        2886 => x"23263101",
        2887 => x"23244101",
        2888 => x"13040600",
        2889 => x"63940502",
        2890 => x"03248101",
        2891 => x"8320c101",
        2892 => x"83244101",
        2893 => x"03290101",
        2894 => x"8329c100",
        2895 => x"032a8100",
        2896 => x"93050600",
        2897 => x"13010102",
        2898 => x"6ff0dfe6",
        2899 => x"63180602",
        2900 => x"eff0dfd6",
        2901 => x"93040000",
        2902 => x"8320c101",
        2903 => x"03248101",
        2904 => x"03290101",
        2905 => x"8329c100",
        2906 => x"032a8100",
        2907 => x"13850400",
        2908 => x"83244101",
        2909 => x"13010102",
        2910 => x"67800000",
        2911 => x"130a0500",
        2912 => x"13890500",
        2913 => x"ef00400a",
        2914 => x"93090500",
        2915 => x"63688500",
        2916 => x"93571500",
        2917 => x"93040900",
        2918 => x"e3e087fc",
        2919 => x"93050400",
        2920 => x"13050a00",
        2921 => x"eff01fe1",
        2922 => x"93040500",
        2923 => x"e30605fa",
        2924 => x"13060400",
        2925 => x"63f48900",
        2926 => x"13860900",
        2927 => x"93050900",
        2928 => x"13850400",
        2929 => x"efe01fae",
        2930 => x"93050900",
        2931 => x"13050a00",
        2932 => x"eff0dfce",
        2933 => x"6ff05ff8",
        2934 => x"130101ff",
        2935 => x"23248100",
        2936 => x"23229100",
        2937 => x"13040500",
        2938 => x"13850500",
        2939 => x"23261100",
        2940 => x"23a20188",
        2941 => x"ef00000c",
        2942 => x"9307f0ff",
        2943 => x"6318f500",
        2944 => x"83a74188",
        2945 => x"63840700",
        2946 => x"2320f400",
        2947 => x"8320c100",
        2948 => x"03248100",
        2949 => x"83244100",
        2950 => x"13010101",
        2951 => x"67800000",
        2952 => x"67800000",
        2953 => x"67800000",
        2954 => x"83a7c5ff",
        2955 => x"1385c7ff",
        2956 => x"63d80700",
        2957 => x"b385a500",
        2958 => x"83a70500",
        2959 => x"3305f500",
        2960 => x"67800000",
        2961 => x"9308d005",
        2962 => x"73000000",
        2963 => x"63520502",
        2964 => x"130101ff",
        2965 => x"23248100",
        2966 => x"13040500",
        2967 => x"23261100",
        2968 => x"33048040",
        2969 => x"efe05fc6",
        2970 => x"23208500",
        2971 => x"6f000000",
        2972 => x"6f000000",
        2973 => x"130101ff",
        2974 => x"23261100",
        2975 => x"23248100",
        2976 => x"9308900a",
        2977 => x"73000000",
        2978 => x"13040500",
        2979 => x"635a0500",
        2980 => x"33048040",
        2981 => x"efe05fc3",
        2982 => x"23208500",
        2983 => x"1304f0ff",
        2984 => x"8320c100",
        2985 => x"13050400",
        2986 => x"03248100",
        2987 => x"13010101",
        2988 => x"67800000",
        2989 => x"83a70189",
        2990 => x"130101ff",
        2991 => x"23261100",
        2992 => x"93060500",
        2993 => x"13870189",
        2994 => x"639c0702",
        2995 => x"9308600d",
        2996 => x"13050000",
        2997 => x"73000000",
        2998 => x"9307f0ff",
        2999 => x"6310f502",
        3000 => x"efe09fbe",
        3001 => x"9307c000",
        3002 => x"2320f500",
        3003 => x"1305f0ff",
        3004 => x"8320c100",
        3005 => x"13010101",
        3006 => x"67800000",
        3007 => x"2320a700",
        3008 => x"83270700",
        3009 => x"9308600d",
        3010 => x"b386f600",
        3011 => x"13850600",
        3012 => x"73000000",
        3013 => x"e316d5fc",
        3014 => x"2320a700",
        3015 => x"13850700",
        3016 => x"6ff01ffd",
        3017 => x"10000000",
        3018 => x"00000000",
        3019 => x"037a5200",
        3020 => x"017c0101",
        3021 => x"1b0d0200",
        3022 => x"10000000",
        3023 => x"18000000",
        3024 => x"88d8ffff",
        3025 => x"78040000",
        3026 => x"00000000",
        3027 => x"10000000",
        3028 => x"00000000",
        3029 => x"037a5200",
        3030 => x"017c0101",
        3031 => x"1b0d0200",
        3032 => x"10000000",
        3033 => x"18000000",
        3034 => x"d8dcffff",
        3035 => x"50040000",
        3036 => x"00000000",
        3037 => x"10000000",
        3038 => x"00000000",
        3039 => x"037a5200",
        3040 => x"017c0101",
        3041 => x"1b0d0200",
        3042 => x"10000000",
        3043 => x"18000000",
        3044 => x"00e1ffff",
        3045 => x"30040000",
        3046 => x"00000000",
        3047 => x"10000000",
        3048 => x"00000000",
        3049 => x"037a5200",
        3050 => x"017c0101",
        3051 => x"1b0d0200",
        3052 => x"10000000",
        3053 => x"18000000",
        3054 => x"08e5ffff",
        3055 => x"e4030000",
        3056 => x"00000000",
        3057 => x"2c020000",
        3058 => x"9c010000",
        3059 => x"9c010000",
        3060 => x"9c010000",
        3061 => x"9c010000",
        3062 => x"10020000",
        3063 => x"9c010000",
        3064 => x"d0010000",
        3065 => x"9c010000",
        3066 => x"9c010000",
        3067 => x"d0010000",
        3068 => x"9c010000",
        3069 => x"9c010000",
        3070 => x"9c010000",
        3071 => x"9c010000",
        3072 => x"9c010000",
        3073 => x"9c010000",
        3074 => x"9c010000",
        3075 => x"80010000",
        3076 => x"40050000",
        3077 => x"28050000",
        3078 => x"28050000",
        3079 => x"28050000",
        3080 => x"28050000",
        3081 => x"58050000",
        3082 => x"ac050000",
        3083 => x"d4050000",
        3084 => x"28050000",
        3085 => x"28050000",
        3086 => x"28050000",
        3087 => x"28050000",
        3088 => x"28050000",
        3089 => x"28050000",
        3090 => x"28050000",
        3091 => x"28050000",
        3092 => x"28050000",
        3093 => x"28050000",
        3094 => x"28050000",
        3095 => x"28050000",
        3096 => x"28050000",
        3097 => x"28050000",
        3098 => x"c8040000",
        3099 => x"c8040000",
        3100 => x"28050000",
        3101 => x"28050000",
        3102 => x"28050000",
        3103 => x"28050000",
        3104 => x"28050000",
        3105 => x"28050000",
        3106 => x"28050000",
        3107 => x"28050000",
        3108 => x"28050000",
        3109 => x"28050000",
        3110 => x"28050000",
        3111 => x"28050000",
        3112 => x"58050000",
        3113 => x"40050000",
        3114 => x"7c050000",
        3115 => x"94050000",
        3116 => x"28050000",
        3117 => x"28050000",
        3118 => x"28050000",
        3119 => x"28050000",
        3120 => x"28050000",
        3121 => x"28050000",
        3122 => x"64050000",
        3123 => x"28050000",
        3124 => x"28050000",
        3125 => x"28050000",
        3126 => x"28050000",
        3127 => x"c8040000",
        3128 => x"c8040000",
        3129 => x"00010202",
        3130 => x"03030303",
        3131 => x"04040404",
        3132 => x"04040404",
        3133 => x"05050505",
        3134 => x"05050505",
        3135 => x"05050505",
        3136 => x"05050505",
        3137 => x"06060606",
        3138 => x"06060606",
        3139 => x"06060606",
        3140 => x"06060606",
        3141 => x"06060606",
        3142 => x"06060606",
        3143 => x"06060606",
        3144 => x"06060606",
        3145 => x"07070707",
        3146 => x"07070707",
        3147 => x"07070707",
        3148 => x"07070707",
        3149 => x"07070707",
        3150 => x"07070707",
        3151 => x"07070707",
        3152 => x"07070707",
        3153 => x"07070707",
        3154 => x"07070707",
        3155 => x"07070707",
        3156 => x"07070707",
        3157 => x"07070707",
        3158 => x"07070707",
        3159 => x"07070707",
        3160 => x"07070707",
        3161 => x"08080808",
        3162 => x"08080808",
        3163 => x"08080808",
        3164 => x"08080808",
        3165 => x"08080808",
        3166 => x"08080808",
        3167 => x"08080808",
        3168 => x"08080808",
        3169 => x"08080808",
        3170 => x"08080808",
        3171 => x"08080808",
        3172 => x"08080808",
        3173 => x"08080808",
        3174 => x"08080808",
        3175 => x"08080808",
        3176 => x"08080808",
        3177 => x"08080808",
        3178 => x"08080808",
        3179 => x"08080808",
        3180 => x"08080808",
        3181 => x"08080808",
        3182 => x"08080808",
        3183 => x"08080808",
        3184 => x"08080808",
        3185 => x"08080808",
        3186 => x"08080808",
        3187 => x"08080808",
        3188 => x"08080808",
        3189 => x"08080808",
        3190 => x"08080808",
        3191 => x"08080808",
        3192 => x"08080808",
        3193 => x"0d0a0d0a",
        3194 => x"44697370",
        3195 => x"6c617969",
        3196 => x"6e672074",
        3197 => x"68652074",
        3198 => x"696d6520",
        3199 => x"70617373",
        3200 => x"65642073",
        3201 => x"696e6365",
        3202 => x"20726573",
        3203 => x"65740d0a",
        3204 => x"0d0a0000",
        3205 => x"2530356c",
        3206 => x"643a2530",
        3207 => x"366c6420",
        3208 => x"20202530",
        3209 => x"326c643a",
        3210 => x"2530326c",
        3211 => x"643a2530",
        3212 => x"326c640d",
        3213 => x"00000000",
        3214 => x"696e7465",
        3215 => x"72727570",
        3216 => x"74000000",
        3217 => x"52495343",
        3218 => x"2d562052",
        3219 => x"56333249",
        3220 => x"4d206261",
        3221 => x"7265206d",
        3222 => x"6574616c",
        3223 => x"2070726f",
        3224 => x"63657373",
        3225 => x"6f720000",
        3226 => x"54686520",
        3227 => x"48616775",
        3228 => x"6520556e",
        3229 => x"69766572",
        3230 => x"73697479",
        3231 => x"206f6620",
        3232 => x"4170706c",
        3233 => x"69656420",
        3234 => x"53636965",
        3235 => x"6e636573",
        3236 => x"00000000",
        3237 => x"44657061",
        3238 => x"72746d65",
        3239 => x"6e74206f",
        3240 => x"6620456c",
        3241 => x"65637472",
        3242 => x"6963616c",
        3243 => x"20456e67",
        3244 => x"696e6565",
        3245 => x"72696e67",
        3246 => x"00000000",
        3247 => x"4a2e452e",
        3248 => x"4a2e206f",
        3249 => x"70206465",
        3250 => x"6e204272",
        3251 => x"6f757700",
        3252 => x"3c627265",
        3253 => x"616b3e0d",
        3254 => x"0a000000",
        3255 => x"0d0a4542",
        3256 => x"5245414b",
        3257 => x"21206d69",
        3258 => x"70203d20",
        3259 => x"00000000",
        3260 => x"232d302b",
        3261 => x"20000000",
        3262 => x"686c4c00",
        3263 => x"65666745",
        3264 => x"46470000",
        3265 => x"30313233",
        3266 => x"34353637",
        3267 => x"38394142",
        3268 => x"43444546",
        3269 => x"00000000",
        3270 => x"30313233",
        3271 => x"34353637",
        3272 => x"38396162",
        3273 => x"63646566",
        3274 => x"00000000",
        3275 => x"e8250000",
        3276 => x"08260000",
        3277 => x"b4250000",
        3278 => x"b4250000",
        3279 => x"b4250000",
        3280 => x"b4250000",
        3281 => x"08260000",
        3282 => x"b4250000",
        3283 => x"b4250000",
        3284 => x"b4250000",
        3285 => x"b4250000",
        3286 => x"f4270000",
        3287 => x"60260000",
        3288 => x"70270000",
        3289 => x"b4250000",
        3290 => x"b4250000",
        3291 => x"3c280000",
        3292 => x"b4250000",
        3293 => x"60260000",
        3294 => x"b4250000",
        3295 => x"b4250000",
        3296 => x"7c270000",
        3297 => x"18000020",
        3298 => x"38320000",
        3299 => x"44320000",
        3300 => x"68320000",
        3301 => x"94320000",
        3302 => x"bc320000",
        3303 => x"00000000",
        3304 => x"00000000",
        3305 => x"00000000",
        3306 => x"00000000",
        3307 => x"00000000",
        3308 => x"00000000",
        3309 => x"00000000",
        3310 => x"00000000",
        3311 => x"00000000",
        3312 => x"00000000",
        3313 => x"00000000",
        3314 => x"00000000",
        3315 => x"00000000",
        3316 => x"00000000",
        3317 => x"00000000",
        3318 => x"00000000",
        3319 => x"00000000",
        3320 => x"00000000",
        3321 => x"00000000",
        3322 => x"00000000",
        3323 => x"00000000",
        3324 => x"00000000",
        3325 => x"00000000",
        3326 => x"00000000",
        3327 => x"00000000",
        3328 => x"80000020",
        3329 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
