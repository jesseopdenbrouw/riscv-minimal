-- srec2vhdl table generator
-- for input file malloc.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17410020",
           3 => x"130181ff",
           4 => x"93804186",
           5 => x"93844187",
           6 => x"b7170000",
           7 => x"13898796",
           8 => x"6f004001",
           9 => x"23a00000",
          10 => x"93870000",
          11 => x"93804700",
          12 => x"83a70700",
          13 => x"e3e890fe",
          14 => x"b7070020",
          15 => x"93800700",
          16 => x"93844186",
          17 => x"6f004001",
          18 => x"83270900",
          19 => x"23a0f000",
          20 => x"93804000",
          21 => x"13094900",
          22 => x"e3e890fe",
          23 => x"13894186",
          24 => x"b7170000",
          25 => x"93804796",
          26 => x"b7170000",
          27 => x"93848796",
          28 => x"6f00c001",
          29 => x"83a70000",
          30 => x"2320f900",
          31 => x"93804000",
          32 => x"93070900",
          33 => x"13894700",
          34 => x"83a70700",
          35 => x"e3e490fe",
          36 => x"ef00002b",
          37 => x"ef00c000",
          38 => x"13050000",
          39 => x"ef004026",
          40 => x"130101fd",
          41 => x"23261102",
          42 => x"23248102",
          43 => x"13040103",
          44 => x"13054006",
          45 => x"ef008032",
          46 => x"93070500",
          47 => x"232ef4fc",
          48 => x"232604fe",
          49 => x"6f004002",
          50 => x"8327c4fe",
          51 => x"0327c4fd",
          52 => x"b307f700",
          53 => x"13071004",
          54 => x"2380e700",
          55 => x"8327c4fe",
          56 => x"93871700",
          57 => x"2326f4fe",
          58 => x"0327c4fe",
          59 => x"93073006",
          60 => x"e3dce7fc",
          61 => x"0325c4fd",
          62 => x"ef00002f",
          63 => x"13052003",
          64 => x"ef00c02d",
          65 => x"93070500",
          66 => x"232ef4fc",
          67 => x"232404fe",
          68 => x"6f000003",
          69 => x"832784fe",
          70 => x"13f7f70f",
          71 => x"832784fe",
          72 => x"8326c4fd",
          73 => x"b387f600",
          74 => x"13071704",
          75 => x"1377f70f",
          76 => x"2380e700",
          77 => x"832784fe",
          78 => x"93871700",
          79 => x"2324f4fe",
          80 => x"032784fe",
          81 => x"93071003",
          82 => x"e3d6e7fc",
          83 => x"0325c4fd",
          84 => x"ef008029",
          85 => x"13054006",
          86 => x"ef004028",
          87 => x"93070500",
          88 => x"232cf4fc",
          89 => x"232204fe",
          90 => x"6f008002",
          91 => x"832744fe",
          92 => x"93972700",
          93 => x"032784fd",
          94 => x"b307f700",
          95 => x"1307f0ff",
          96 => x"23a0e700",
          97 => x"832744fe",
          98 => x"93871700",
          99 => x"2322f4fe",
         100 => x"032744fe",
         101 => x"93072006",
         102 => x"e3dae7fc",
         103 => x"032584fd",
         104 => x"ef008024",
         105 => x"93054000",
         106 => x"13059001",
         107 => x"ef00c013",
         108 => x"93070500",
         109 => x"232af4fc",
         110 => x"232004fe",
         111 => x"6f00c002",
         112 => x"832704fe",
         113 => x"93972700",
         114 => x"032744fd",
         115 => x"b307f700",
         116 => x"37171111",
         117 => x"13071711",
         118 => x"23a0e700",
         119 => x"832704fe",
         120 => x"93871700",
         121 => x"2320f4fe",
         122 => x"032704fe",
         123 => x"93078001",
         124 => x"e3d8e7fc",
         125 => x"93070000",
         126 => x"13850700",
         127 => x"8320c102",
         128 => x"03248102",
         129 => x"13010103",
         130 => x"67800000",
         131 => x"130101fd",
         132 => x"23261102",
         133 => x"23248102",
         134 => x"13040103",
         135 => x"232ea4fc",
         136 => x"b7470020",
         137 => x"13870700",
         138 => x"93070040",
         139 => x"b307f740",
         140 => x"2326f4fe",
         141 => x"8327c4fe",
         142 => x"2324f4fe",
         143 => x"83a70187",
         144 => x"63960700",
         145 => x"13878187",
         146 => x"23a8e186",
         147 => x"03a70187",
         148 => x"8327c4fd",
         149 => x"b307f700",
         150 => x"032784fe",
         151 => x"637ef700",
         152 => x"ef008009",
         153 => x"13070500",
         154 => x"9307c000",
         155 => x"2320f700",
         156 => x"9307f0ff",
         157 => x"6f000002",
         158 => x"83a70187",
         159 => x"2322f4fe",
         160 => x"03a70187",
         161 => x"8327c4fd",
         162 => x"3307f700",
         163 => x"23a8e186",
         164 => x"832744fe",
         165 => x"13850700",
         166 => x"8320c102",
         167 => x"03248102",
         168 => x"13010103",
         169 => x"67800000",
         170 => x"13030500",
         171 => x"630a0600",
         172 => x"2300b300",
         173 => x"1306f6ff",
         174 => x"13031300",
         175 => x"e31a06fe",
         176 => x"67800000",
         177 => x"13060500",
         178 => x"13050000",
         179 => x"93f61500",
         180 => x"63840600",
         181 => x"3305c500",
         182 => x"93d51500",
         183 => x"13161600",
         184 => x"e39605fe",
         185 => x"67800000",
         186 => x"13860500",
         187 => x"93050500",
         188 => x"03a50186",
         189 => x"6f000010",
         190 => x"03a50186",
         191 => x"67800000",
         192 => x"130101ff",
         193 => x"23248100",
         194 => x"23261100",
         195 => x"93070000",
         196 => x"13040500",
         197 => x"63880700",
         198 => x"93050000",
         199 => x"97000000",
         200 => x"e7000000",
         201 => x"b7170000",
         202 => x"03a54796",
         203 => x"83278502",
         204 => x"63840700",
         205 => x"e7800700",
         206 => x"13050400",
         207 => x"ef00805f",
         208 => x"130101ff",
         209 => x"23248100",
         210 => x"23229100",
         211 => x"37140000",
         212 => x"b7140000",
         213 => x"93878496",
         214 => x"13048496",
         215 => x"3304f440",
         216 => x"23202101",
         217 => x"23261100",
         218 => x"13542440",
         219 => x"93848496",
         220 => x"13090000",
         221 => x"63108904",
         222 => x"b7140000",
         223 => x"37140000",
         224 => x"93878496",
         225 => x"13048496",
         226 => x"3304f440",
         227 => x"13542440",
         228 => x"93848496",
         229 => x"13090000",
         230 => x"63188902",
         231 => x"8320c100",
         232 => x"03248100",
         233 => x"83244100",
         234 => x"03290100",
         235 => x"13010101",
         236 => x"67800000",
         237 => x"83a70400",
         238 => x"13091900",
         239 => x"93844400",
         240 => x"e7800700",
         241 => x"6ff01ffb",
         242 => x"83a70400",
         243 => x"13091900",
         244 => x"93844400",
         245 => x"e7800700",
         246 => x"6ff01ffc",
         247 => x"93050500",
         248 => x"03a50186",
         249 => x"6f008020",
         250 => x"93050500",
         251 => x"03a50186",
         252 => x"6f004010",
         253 => x"130101fd",
         254 => x"23229102",
         255 => x"23202103",
         256 => x"23261102",
         257 => x"23248102",
         258 => x"232e3101",
         259 => x"13d90501",
         260 => x"93040500",
         261 => x"93560601",
         262 => x"13850500",
         263 => x"6310090a",
         264 => x"63920604",
         265 => x"93150601",
         266 => x"13150501",
         267 => x"93d50501",
         268 => x"13550501",
         269 => x"eff01fe9",
         270 => x"13060500",
         271 => x"93050600",
         272 => x"13850400",
         273 => x"2326c100",
         274 => x"ef00401a",
         275 => x"13040500",
         276 => x"63020508",
         277 => x"0326c100",
         278 => x"93050000",
         279 => x"eff0dfe4",
         280 => x"6f004007",
         281 => x"13890600",
         282 => x"93890500",
         283 => x"93150601",
         284 => x"13150501",
         285 => x"93d50501",
         286 => x"13550501",
         287 => x"eff09fe4",
         288 => x"13040500",
         289 => x"93150901",
         290 => x"13950901",
         291 => x"93d50501",
         292 => x"13550501",
         293 => x"eff01fe3",
         294 => x"93570401",
         295 => x"3306f500",
         296 => x"93570601",
         297 => x"63920702",
         298 => x"13140401",
         299 => x"13160601",
         300 => x"13540401",
         301 => x"33668600",
         302 => x"6ff05ff8",
         303 => x"63960600",
         304 => x"93090600",
         305 => x"6ff09ffa",
         306 => x"9307c000",
         307 => x"23a0f400",
         308 => x"13040000",
         309 => x"8320c102",
         310 => x"13050400",
         311 => x"03248102",
         312 => x"83244102",
         313 => x"03290102",
         314 => x"8329c101",
         315 => x"13010103",
         316 => x"67800000",
         317 => x"638a050e",
         318 => x"83a7c5ff",
         319 => x"130101fe",
         320 => x"232c8100",
         321 => x"232e1100",
         322 => x"1384c5ff",
         323 => x"63d40700",
         324 => x"3304f400",
         325 => x"2326a100",
         326 => x"ef00c026",
         327 => x"83a74186",
         328 => x"0325c100",
         329 => x"639e0700",
         330 => x"23220400",
         331 => x"23a28186",
         332 => x"03248101",
         333 => x"8320c101",
         334 => x"13010102",
         335 => x"6f00c024",
         336 => x"6374f402",
         337 => x"03260400",
         338 => x"b306c400",
         339 => x"639ad700",
         340 => x"83a60700",
         341 => x"83a74700",
         342 => x"b386c600",
         343 => x"2320d400",
         344 => x"2322f400",
         345 => x"6ff09ffc",
         346 => x"13870700",
         347 => x"83a74700",
         348 => x"63840700",
         349 => x"e37af4fe",
         350 => x"83260700",
         351 => x"3306d700",
         352 => x"63188602",
         353 => x"03260400",
         354 => x"b386c600",
         355 => x"2320d700",
         356 => x"3306d700",
         357 => x"e39ec7f8",
         358 => x"03a60700",
         359 => x"83a74700",
         360 => x"b306d600",
         361 => x"2320d700",
         362 => x"2322f700",
         363 => x"6ff05ff8",
         364 => x"6378c400",
         365 => x"9307c000",
         366 => x"2320f500",
         367 => x"6ff05ff7",
         368 => x"03260400",
         369 => x"b306c400",
         370 => x"639ad700",
         371 => x"83a60700",
         372 => x"83a74700",
         373 => x"b386c600",
         374 => x"2320d400",
         375 => x"2322f400",
         376 => x"23228700",
         377 => x"6ff0dff4",
         378 => x"67800000",
         379 => x"130101fe",
         380 => x"232a9100",
         381 => x"93843500",
         382 => x"93f4c4ff",
         383 => x"23282101",
         384 => x"232e1100",
         385 => x"232c8100",
         386 => x"23263101",
         387 => x"93848400",
         388 => x"9307c000",
         389 => x"13090500",
         390 => x"63f4f406",
         391 => x"9304c000",
         392 => x"63e2b406",
         393 => x"13050900",
         394 => x"ef00c015",
         395 => x"03a74186",
         396 => x"93864186",
         397 => x"13040700",
         398 => x"631a0406",
         399 => x"13848186",
         400 => x"83270400",
         401 => x"639a0700",
         402 => x"93050000",
         403 => x"13050900",
         404 => x"ef00c00e",
         405 => x"2320a400",
         406 => x"93850400",
         407 => x"13050900",
         408 => x"ef00c00d",
         409 => x"9309f0ff",
         410 => x"631a350b",
         411 => x"9307c000",
         412 => x"2320f900",
         413 => x"13050900",
         414 => x"ef000011",
         415 => x"6f000001",
         416 => x"e3d004fa",
         417 => x"9307c000",
         418 => x"2320f900",
         419 => x"13050000",
         420 => x"8320c101",
         421 => x"03248101",
         422 => x"83244101",
         423 => x"03290101",
         424 => x"8329c100",
         425 => x"13010102",
         426 => x"67800000",
         427 => x"83270400",
         428 => x"b3879740",
         429 => x"63ce0704",
         430 => x"1306b000",
         431 => x"637af600",
         432 => x"2320f400",
         433 => x"3304f400",
         434 => x"23209400",
         435 => x"6f000001",
         436 => x"83274400",
         437 => x"631a8702",
         438 => x"23a0f600",
         439 => x"13050900",
         440 => x"ef00800a",
         441 => x"1305b400",
         442 => x"93074400",
         443 => x"137585ff",
         444 => x"3307f540",
         445 => x"e30ef5f8",
         446 => x"3304e400",
         447 => x"b387a740",
         448 => x"2320f400",
         449 => x"6ff0dff8",
         450 => x"2322f700",
         451 => x"6ff01ffd",
         452 => x"13070400",
         453 => x"03244400",
         454 => x"6ff01ff2",
         455 => x"13043500",
         456 => x"1374c4ff",
         457 => x"e30285fa",
         458 => x"b305a440",
         459 => x"13050900",
         460 => x"ef00c000",
         461 => x"e31a35f9",
         462 => x"6ff05ff3",
         463 => x"130101ff",
         464 => x"23248100",
         465 => x"23229100",
         466 => x"13040500",
         467 => x"13850500",
         468 => x"23261100",
         469 => x"23a60186",
         470 => x"eff05fab",
         471 => x"9307f0ff",
         472 => x"6318f500",
         473 => x"83a7c186",
         474 => x"63840700",
         475 => x"2320f400",
         476 => x"8320c100",
         477 => x"03248100",
         478 => x"83244100",
         479 => x"13010101",
         480 => x"67800000",
         481 => x"67800000",
         482 => x"67800000",
         483 => x"130101ff",
         484 => x"23248100",
         485 => x"13840500",
         486 => x"83a50500",
         487 => x"23229100",
         488 => x"23261100",
         489 => x"93040500",
         490 => x"63840500",
         491 => x"eff01ffe",
         492 => x"93050400",
         493 => x"03248100",
         494 => x"8320c100",
         495 => x"13850400",
         496 => x"83244100",
         497 => x"13010101",
         498 => x"6ff0dfd2",
         499 => x"83a70186",
         500 => x"6380a716",
         501 => x"83274502",
         502 => x"130101fe",
         503 => x"232c8100",
         504 => x"232e1100",
         505 => x"232a9100",
         506 => x"23282101",
         507 => x"23263101",
         508 => x"13040500",
         509 => x"63840702",
         510 => x"83a7c700",
         511 => x"93040000",
         512 => x"13090008",
         513 => x"6392070e",
         514 => x"83274402",
         515 => x"83a50700",
         516 => x"63860500",
         517 => x"13050400",
         518 => x"eff0dfcd",
         519 => x"83254401",
         520 => x"63860500",
         521 => x"13050400",
         522 => x"eff0dfcc",
         523 => x"83254402",
         524 => x"63860500",
         525 => x"13050400",
         526 => x"eff0dfcb",
         527 => x"83258403",
         528 => x"63860500",
         529 => x"13050400",
         530 => x"eff0dfca",
         531 => x"8325c403",
         532 => x"63860500",
         533 => x"13050400",
         534 => x"eff0dfc9",
         535 => x"83250404",
         536 => x"63860500",
         537 => x"13050400",
         538 => x"eff0dfc8",
         539 => x"8325c405",
         540 => x"63860500",
         541 => x"13050400",
         542 => x"eff0dfc7",
         543 => x"83258405",
         544 => x"63860500",
         545 => x"13050400",
         546 => x"eff0dfc6",
         547 => x"83254403",
         548 => x"63860500",
         549 => x"13050400",
         550 => x"eff0dfc5",
         551 => x"83278401",
         552 => x"638a0706",
         553 => x"83278402",
         554 => x"13050400",
         555 => x"e7800700",
         556 => x"83258404",
         557 => x"63800506",
         558 => x"13050400",
         559 => x"03248101",
         560 => x"8320c101",
         561 => x"83244101",
         562 => x"03290101",
         563 => x"8329c100",
         564 => x"13010102",
         565 => x"6ff09feb",
         566 => x"b3859500",
         567 => x"83a50500",
         568 => x"63900502",
         569 => x"93844400",
         570 => x"83274402",
         571 => x"83a5c700",
         572 => x"e39424ff",
         573 => x"13050400",
         574 => x"eff0dfbf",
         575 => x"6ff0dff0",
         576 => x"83a90500",
         577 => x"13050400",
         578 => x"eff0dfbe",
         579 => x"93850900",
         580 => x"6ff01ffd",
         581 => x"8320c101",
         582 => x"03248101",
         583 => x"83244101",
         584 => x"03290101",
         585 => x"8329c100",
         586 => x"13010102",
         587 => x"67800000",
         588 => x"67800000",
         589 => x"9308d005",
         590 => x"73000000",
         591 => x"63520502",
         592 => x"130101ff",
         593 => x"23248100",
         594 => x"13040500",
         595 => x"23261100",
         596 => x"33048040",
         597 => x"eff05f9a",
         598 => x"23208500",
         599 => x"6f000000",
         600 => x"6f000000",
         601 => x"00000020",
         602 => x"00000000",
         603 => x"00000000",
         604 => x"00000000",
         605 => x"00000000",
         606 => x"00000000",
         607 => x"00000000",
         608 => x"00000000",
         609 => x"00000000",
         610 => x"00000000",
         611 => x"00000000",
         612 => x"00000000",
         613 => x"00000000",
         614 => x"00000000",
         615 => x"00000000",
         616 => x"00000000",
         617 => x"00000000",
         618 => x"00000000",
         619 => x"00000000",
         620 => x"00000000",
         621 => x"00000000",
         622 => x"00000000",
         623 => x"00000000",
         624 => x"00000000",
         625 => x"00000000",
         626 => x"00000020",
        others => (others => '-')
    );
end package processor_common_rom;
