-- srec2vhdl table generator
-- for input file float.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17410020",
           3 => x"130181ff",
           4 => x"93864186",
           5 => x"13874186",
           6 => x"63f8e602",
           7 => x"1307f7ff",
           8 => x"3307d740",
           9 => x"1377c7ff",
          10 => x"13074700",
          11 => x"b386e600",
          12 => x"93874186",
          13 => x"23a00700",
          14 => x"13870700",
          15 => x"03270700",
          16 => x"93874700",
          17 => x"e398d7fe",
          18 => x"37070020",
          19 => x"93050700",
          20 => x"93874186",
          21 => x"63fcf502",
          22 => x"9386f7ff",
          23 => x"b386b640",
          24 => x"93f6c6ff",
          25 => x"93864600",
          26 => x"b385d500",
          27 => x"b7160000",
          28 => x"93864602",
          29 => x"13070700",
          30 => x"03a60600",
          31 => x"13074700",
          32 => x"93864600",
          33 => x"232ec7fe",
          34 => x"e318b7fe",
          35 => x"37170000",
          36 => x"b7160000",
          37 => x"930547ed",
          38 => x"93864602",
          39 => x"63fcd502",
          40 => x"9386f6ff",
          41 => x"b386b640",
          42 => x"93f6c6ff",
          43 => x"93864600",
          44 => x"b385d500",
          45 => x"130747ed",
          46 => x"03260700",
          47 => x"93860700",
          48 => x"13074700",
          49 => x"23a0c700",
          50 => x"83a60600",
          51 => x"93874700",
          52 => x"e394e5fe",
          53 => x"ef00d052",
          54 => x"ef009048",
          55 => x"13050000",
          56 => x"ef00104e",
          57 => x"37078000",
          58 => x"130101ff",
          59 => x"1307f7ff",
          60 => x"b377a700",
          61 => x"23248100",
          62 => x"23229100",
          63 => x"13547501",
          64 => x"9354f501",
          65 => x"13d57501",
          66 => x"3377b700",
          67 => x"1374f40f",
          68 => x"1375f50f",
          69 => x"23261100",
          70 => x"23202101",
          71 => x"93d5f501",
          72 => x"93973700",
          73 => x"13173700",
          74 => x"b306a440",
          75 => x"6396b418",
          76 => x"6358d00a",
          77 => x"63100504",
          78 => x"63000702",
          79 => x"9306f4ff",
          80 => x"63980600",
          81 => x"b387e700",
          82 => x"13041000",
          83 => x"6f000006",
          84 => x"1306f00f",
          85 => x"6318c402",
          86 => x"13f77700",
          87 => x"630a0734",
          88 => x"13f7f700",
          89 => x"93064000",
          90 => x"6304d734",
          91 => x"93874700",
          92 => x"6f000034",
          93 => x"1306f00f",
          94 => x"e300c4fe",
          95 => x"37060004",
          96 => x"3367c700",
          97 => x"9305b001",
          98 => x"13061000",
          99 => x"63ced500",
         100 => x"13060002",
         101 => x"b355d700",
         102 => x"b306d640",
         103 => x"3317d700",
         104 => x"3337e000",
         105 => x"33e6e500",
         106 => x"b387c700",
         107 => x"37070004",
         108 => x"33f7e700",
         109 => x"e30207fa",
         110 => x"13041400",
         111 => x"1307f00f",
         112 => x"6306e42e",
         113 => x"3707007e",
         114 => x"93f61700",
         115 => x"1307f7ff",
         116 => x"93d71700",
         117 => x"b3f7e700",
         118 => x"b3e7d700",
         119 => x"6ff0dff7",
         120 => x"63860606",
         121 => x"b3068540",
         122 => x"63100402",
         123 => x"6386072a",
         124 => x"1386f6ff",
         125 => x"e30806f4",
         126 => x"9305f00f",
         127 => x"6390b602",
         128 => x"93070700",
         129 => x"6f000021",
         130 => x"1306f00f",
         131 => x"e30ac5fe",
         132 => x"37060004",
         133 => x"b3e7c700",
         134 => x"13860600",
         135 => x"9305b001",
         136 => x"93061000",
         137 => x"63cec500",
         138 => x"93060002",
         139 => x"b386c640",
         140 => x"b3d5c700",
         141 => x"b397d700",
         142 => x"b337f000",
         143 => x"b3e6f500",
         144 => x"b387e600",
         145 => x"13040500",
         146 => x"6ff05ff6",
         147 => x"93061400",
         148 => x"13f6e60f",
         149 => x"63160604",
         150 => x"63180402",
         151 => x"63820724",
         152 => x"e30c07ee",
         153 => x"b387e700",
         154 => x"37070004",
         155 => x"33f7e700",
         156 => x"e30407ee",
         157 => x"370700fc",
         158 => x"1307f7ff",
         159 => x"b3f7e700",
         160 => x"13041000",
         161 => x"6ff05fed",
         162 => x"e38c07f6",
         163 => x"63040718",
         164 => x"93040000",
         165 => x"b7070002",
         166 => x"1304f00f",
         167 => x"6f004021",
         168 => x"1306f00f",
         169 => x"6382c620",
         170 => x"3387e700",
         171 => x"93571700",
         172 => x"13840600",
         173 => x"6ff05fea",
         174 => x"635ed006",
         175 => x"63120506",
         176 => x"e30c07e8",
         177 => x"9306f4ff",
         178 => x"63980600",
         179 => x"b387e740",
         180 => x"13041000",
         181 => x"6f004003",
         182 => x"1306f00f",
         183 => x"e30ec4e6",
         184 => x"9305b001",
         185 => x"13061000",
         186 => x"63ced500",
         187 => x"13060002",
         188 => x"b355d700",
         189 => x"b306d640",
         190 => x"3317d700",
         191 => x"3337e000",
         192 => x"33e6e500",
         193 => x"b387c740",
         194 => x"37090004",
         195 => x"33f72701",
         196 => x"e30407e4",
         197 => x"1309f9ff",
         198 => x"33f92701",
         199 => x"6f008011",
         200 => x"1306f00f",
         201 => x"e30ac4e2",
         202 => x"37060004",
         203 => x"3367c700",
         204 => x"6ff01ffb",
         205 => x"63800608",
         206 => x"b3068540",
         207 => x"63180402",
         208 => x"6382071e",
         209 => x"1386f6ff",
         210 => x"63180600",
         211 => x"b307f740",
         212 => x"93840500",
         213 => x"6ff0dff7",
         214 => x"1308f00f",
         215 => x"63920603",
         216 => x"93070700",
         217 => x"1304f00f",
         218 => x"6f00c006",
         219 => x"1306f00f",
         220 => x"e308c5fe",
         221 => x"37060004",
         222 => x"b3e7c700",
         223 => x"13860600",
         224 => x"1308b001",
         225 => x"93061000",
         226 => x"634ec800",
         227 => x"93060002",
         228 => x"b386c640",
         229 => x"33d8c700",
         230 => x"b397d700",
         231 => x"b337f000",
         232 => x"b366f800",
         233 => x"b307d740",
         234 => x"13040500",
         235 => x"93840500",
         236 => x"6ff09ff5",
         237 => x"93061400",
         238 => x"93f6e60f",
         239 => x"63900606",
         240 => x"63120404",
         241 => x"639c0700",
         242 => x"93040000",
         243 => x"6302070e",
         244 => x"93070700",
         245 => x"93840500",
         246 => x"6ff01fd8",
         247 => x"e30e07d6",
         248 => x"b386e740",
         249 => x"37060004",
         250 => x"33f6c600",
         251 => x"b307f740",
         252 => x"e31206fe",
         253 => x"93070000",
         254 => x"63820608",
         255 => x"93870600",
         256 => x"6ff09fd5",
         257 => x"e39407e8",
         258 => x"e30407e8",
         259 => x"93070700",
         260 => x"93840500",
         261 => x"1304f00f",
         262 => x"6ff01fd4",
         263 => x"3389e740",
         264 => x"b7060004",
         265 => x"b376d900",
         266 => x"63840604",
         267 => x"3309f740",
         268 => x"93840500",
         269 => x"13050900",
         270 => x"ef00d00d",
         271 => x"1305b5ff",
         272 => x"3319a900",
         273 => x"63408504",
         274 => x"33058540",
         275 => x"13051500",
         276 => x"13070002",
         277 => x"3307a740",
         278 => x"b357a900",
         279 => x"3319e900",
         280 => x"33392001",
         281 => x"b3e72701",
         282 => x"13040000",
         283 => x"6ff0dfce",
         284 => x"e31209fc",
         285 => x"93070000",
         286 => x"13040000",
         287 => x"93040000",
         288 => x"6f000003",
         289 => x"b70700fc",
         290 => x"9387f7ff",
         291 => x"3304a440",
         292 => x"b377f900",
         293 => x"6ff05fcc",
         294 => x"93070700",
         295 => x"6ff05fe1",
         296 => x"93070700",
         297 => x"6ff05fcb",
         298 => x"1304f00f",
         299 => x"93070000",
         300 => x"37070004",
         301 => x"33f7e700",
         302 => x"630e0700",
         303 => x"13041400",
         304 => x"1307f00f",
         305 => x"6306e406",
         306 => x"370700fc",
         307 => x"1307f7ff",
         308 => x"b3f7e700",
         309 => x"1307f00f",
         310 => x"93d73700",
         311 => x"6318e400",
         312 => x"63860700",
         313 => x"b7074000",
         314 => x"93040000",
         315 => x"13147401",
         316 => x"3707807f",
         317 => x"93979700",
         318 => x"3374e400",
         319 => x"93d79700",
         320 => x"3364f400",
         321 => x"1395f401",
         322 => x"8320c100",
         323 => x"3365a400",
         324 => x"03248100",
         325 => x"83244100",
         326 => x"03290100",
         327 => x"13010101",
         328 => x"67800000",
         329 => x"93070700",
         330 => x"13840600",
         331 => x"6ff09fea",
         332 => x"93070000",
         333 => x"6ff01ffa",
         334 => x"130101fd",
         335 => x"23229102",
         336 => x"93547501",
         337 => x"232e3101",
         338 => x"232a5101",
         339 => x"23286101",
         340 => x"931a9500",
         341 => x"23261102",
         342 => x"23248102",
         343 => x"23202103",
         344 => x"232c4101",
         345 => x"23267101",
         346 => x"23248101",
         347 => x"93f4f40f",
         348 => x"138b0500",
         349 => x"93da9a00",
         350 => x"9359f501",
         351 => x"63840408",
         352 => x"9307f00f",
         353 => x"6380f40a",
         354 => x"939a3a00",
         355 => x"b7070004",
         356 => x"b3eafa00",
         357 => x"938414f8",
         358 => x"930b0000",
         359 => x"93577b01",
         360 => x"13149b00",
         361 => x"93f7f70f",
         362 => x"13549400",
         363 => x"135bfb01",
         364 => x"638a0708",
         365 => x"1307f00f",
         366 => x"6386e70a",
         367 => x"13143400",
         368 => x"37070004",
         369 => x"3364e400",
         370 => x"938717f8",
         371 => x"13070000",
         372 => x"338af440",
         373 => x"93972b00",
         374 => x"b3e7e700",
         375 => x"9387f7ff",
         376 => x"9306e000",
         377 => x"33c96901",
         378 => x"63eef608",
         379 => x"b7160000",
         380 => x"93972700",
         381 => x"938646ed",
         382 => x"b387d700",
         383 => x"83a70700",
         384 => x"67800700",
         385 => x"638a0a02",
         386 => x"13850a00",
         387 => x"ef008070",
         388 => x"9307b5ff",
         389 => x"9304a0f8",
         390 => x"b39afa00",
         391 => x"b384a440",
         392 => x"6ff09ff7",
         393 => x"9304f00f",
         394 => x"930b2000",
         395 => x"e3880af6",
         396 => x"930b3000",
         397 => x"6ff09ff6",
         398 => x"93040000",
         399 => x"930b1000",
         400 => x"6ff0dff5",
         401 => x"630a0402",
         402 => x"13050400",
         403 => x"ef00806c",
         404 => x"9307b5ff",
         405 => x"3314f400",
         406 => x"9307a0f8",
         407 => x"b387a740",
         408 => x"6ff0dff6",
         409 => x"9307f00f",
         410 => x"13072000",
         411 => x"e30204f6",
         412 => x"13073000",
         413 => x"6ff0dff5",
         414 => x"93070000",
         415 => x"13071000",
         416 => x"6ff01ff5",
         417 => x"131c5400",
         418 => x"63fa8a16",
         419 => x"130afaff",
         420 => x"13040000",
         421 => x"135b0c01",
         422 => x"b7090100",
         423 => x"93050b00",
         424 => x"9389f9ff",
         425 => x"13850a00",
         426 => x"ef00005c",
         427 => x"b3793c01",
         428 => x"93050500",
         429 => x"930b0500",
         430 => x"13850900",
         431 => x"ef000058",
         432 => x"93040500",
         433 => x"93050b00",
         434 => x"13850a00",
         435 => x"ef00405e",
         436 => x"93570401",
         437 => x"13150501",
         438 => x"b3e7a700",
         439 => x"13840b00",
         440 => x"63fe9700",
         441 => x"b3878701",
         442 => x"1384fbff",
         443 => x"63e88701",
         444 => x"63f69700",
         445 => x"1384ebff",
         446 => x"b3878701",
         447 => x"b3849740",
         448 => x"93050b00",
         449 => x"13850400",
         450 => x"ef000056",
         451 => x"93050500",
         452 => x"930a0500",
         453 => x"13850900",
         454 => x"ef004052",
         455 => x"93090500",
         456 => x"93050b00",
         457 => x"13850400",
         458 => x"ef008058",
         459 => x"93170501",
         460 => x"13870a00",
         461 => x"63fe3701",
         462 => x"b3878701",
         463 => x"1387faff",
         464 => x"63e88701",
         465 => x"63f63701",
         466 => x"1387eaff",
         467 => x"b3878701",
         468 => x"13140401",
         469 => x"b3873741",
         470 => x"3364e400",
         471 => x"b337f000",
         472 => x"3364f400",
         473 => x"1307fa07",
         474 => x"6354e00e",
         475 => x"93777400",
         476 => x"638a0700",
         477 => x"9377f400",
         478 => x"93064000",
         479 => x"6384d700",
         480 => x"13044400",
         481 => x"b7070008",
         482 => x"b377f400",
         483 => x"638a0700",
         484 => x"b70700f8",
         485 => x"9387f7ff",
         486 => x"3374f400",
         487 => x"13070a08",
         488 => x"9307e00f",
         489 => x"63c4e708",
         490 => x"93573400",
         491 => x"8320c102",
         492 => x"03248102",
         493 => x"13177701",
         494 => x"b706807f",
         495 => x"93979700",
         496 => x"3377d700",
         497 => x"93d79700",
         498 => x"1315f901",
         499 => x"3367f700",
         500 => x"83244102",
         501 => x"03290102",
         502 => x"8329c101",
         503 => x"032a8101",
         504 => x"832a4101",
         505 => x"032b0101",
         506 => x"832bc100",
         507 => x"032c8100",
         508 => x"3365a700",
         509 => x"13010103",
         510 => x"67800000",
         511 => x"1394fa01",
         512 => x"93da1a00",
         513 => x"6ff01fe9",
         514 => x"13890900",
         515 => x"13840a00",
         516 => x"13870b00",
         517 => x"93073000",
         518 => x"6308f708",
         519 => x"93071000",
         520 => x"630cf708",
         521 => x"93072000",
         522 => x"e31ef7f2",
         523 => x"93070000",
         524 => x"1307f00f",
         525 => x"6ff09ff7",
         526 => x"13090b00",
         527 => x"6ff09ffd",
         528 => x"37044000",
         529 => x"13090000",
         530 => x"13073000",
         531 => x"6ff09ffc",
         532 => x"93071000",
         533 => x"b387e740",
         534 => x"1307b001",
         535 => x"634ef704",
         536 => x"9304ea09",
         537 => x"b357f400",
         538 => x"33149400",
         539 => x"33348000",
         540 => x"b3e78700",
         541 => x"13f77700",
         542 => x"630a0700",
         543 => x"13f7f700",
         544 => x"93064000",
         545 => x"6304d700",
         546 => x"93874700",
         547 => x"37070004",
         548 => x"33f7e700",
         549 => x"93d73700",
         550 => x"e30a07f0",
         551 => x"93070000",
         552 => x"13071000",
         553 => x"6ff09ff0",
         554 => x"b7074000",
         555 => x"1307f00f",
         556 => x"13090000",
         557 => x"6ff09fef",
         558 => x"93070000",
         559 => x"13070000",
         560 => x"6ff0dfee",
         561 => x"130101fe",
         562 => x"23282101",
         563 => x"13597501",
         564 => x"232a9100",
         565 => x"23263101",
         566 => x"23225101",
         567 => x"93149500",
         568 => x"232e1100",
         569 => x"232c8100",
         570 => x"23244101",
         571 => x"1379f90f",
         572 => x"938a0500",
         573 => x"93d49400",
         574 => x"9359f501",
         575 => x"6302091c",
         576 => x"9307f00f",
         577 => x"630ef91c",
         578 => x"93943400",
         579 => x"b7070004",
         580 => x"b3e4f400",
         581 => x"130919f8",
         582 => x"130a0000",
         583 => x"93d77a01",
         584 => x"13949a00",
         585 => x"93f7f70f",
         586 => x"13549400",
         587 => x"93dafa01",
         588 => x"6388071c",
         589 => x"1307f00f",
         590 => x"6384e71e",
         591 => x"13143400",
         592 => x"37070004",
         593 => x"3364e400",
         594 => x"938717f8",
         595 => x"93060000",
         596 => x"3309f900",
         597 => x"93172a00",
         598 => x"b3e7d700",
         599 => x"1307a000",
         600 => x"33c85901",
         601 => x"93081900",
         602 => x"6344f722",
         603 => x"13072000",
         604 => x"6348f71c",
         605 => x"9387f7ff",
         606 => x"13071000",
         607 => x"6374f71e",
         608 => x"b70e0100",
         609 => x"1383feff",
         610 => x"93df0401",
         611 => x"135f0401",
         612 => x"b3f46400",
         613 => x"33746400",
         614 => x"13850400",
         615 => x"93050400",
         616 => x"ef00c029",
         617 => x"13070500",
         618 => x"93050f00",
         619 => x"13850400",
         620 => x"ef00c028",
         621 => x"93070500",
         622 => x"93050400",
         623 => x"13850f00",
         624 => x"ef00c027",
         625 => x"130e0500",
         626 => x"93050f00",
         627 => x"13850f00",
         628 => x"ef00c026",
         629 => x"13540701",
         630 => x"b387c701",
         631 => x"3304f400",
         632 => x"93060500",
         633 => x"6374c401",
         634 => x"b306d501",
         635 => x"b3776400",
         636 => x"33776700",
         637 => x"93970701",
         638 => x"b387e700",
         639 => x"13976700",
         640 => x"13540401",
         641 => x"3337e000",
         642 => x"93d7a701",
         643 => x"3304d400",
         644 => x"b367f700",
         645 => x"13146400",
         646 => x"3364f400",
         647 => x"b7070008",
         648 => x"b377f400",
         649 => x"638e0718",
         650 => x"93571400",
         651 => x"13741400",
         652 => x"33e48700",
         653 => x"1387f807",
         654 => x"6358e018",
         655 => x"93777400",
         656 => x"638a0700",
         657 => x"9377f400",
         658 => x"93064000",
         659 => x"6384d700",
         660 => x"13044400",
         661 => x"b7070008",
         662 => x"b377f400",
         663 => x"638a0700",
         664 => x"b70700f8",
         665 => x"9387f7ff",
         666 => x"3374f400",
         667 => x"13870808",
         668 => x"9307e00f",
         669 => x"63cee71a",
         670 => x"93573400",
         671 => x"8320c101",
         672 => x"03248101",
         673 => x"13177701",
         674 => x"b706807f",
         675 => x"93979700",
         676 => x"3377d700",
         677 => x"93d79700",
         678 => x"3367f700",
         679 => x"1315f801",
         680 => x"83244101",
         681 => x"03290101",
         682 => x"8329c100",
         683 => x"032a8100",
         684 => x"832a4100",
         685 => x"3365a700",
         686 => x"13010102",
         687 => x"67800000",
         688 => x"638a0402",
         689 => x"13850400",
         690 => x"ef00c024",
         691 => x"9307b5ff",
         692 => x"1309a0f8",
         693 => x"b394f400",
         694 => x"3309a940",
         695 => x"6ff0dfe3",
         696 => x"1309f00f",
         697 => x"130a2000",
         698 => x"e38a04e2",
         699 => x"130a3000",
         700 => x"6ff0dfe2",
         701 => x"13090000",
         702 => x"130a1000",
         703 => x"6ff01fe2",
         704 => x"630a0402",
         705 => x"13050400",
         706 => x"ef00c020",
         707 => x"9307b5ff",
         708 => x"3314f400",
         709 => x"9307a0f8",
         710 => x"b387a740",
         711 => x"6ff01fe3",
         712 => x"9307f00f",
         713 => x"93062000",
         714 => x"e30404e2",
         715 => x"93063000",
         716 => x"6ff01fe2",
         717 => x"93070000",
         718 => x"93061000",
         719 => x"6ff05fe1",
         720 => x"13071000",
         721 => x"b317f700",
         722 => x"13f70753",
         723 => x"631c0704",
         724 => x"13f70724",
         725 => x"6316070c",
         726 => x"93f78708",
         727 => x"e38207e2",
         728 => x"13880a00",
         729 => x"13062000",
         730 => x"93070000",
         731 => x"1307f00f",
         732 => x"e386c6f0",
         733 => x"93073000",
         734 => x"6384f60a",
         735 => x"93071000",
         736 => x"e39af6ea",
         737 => x"93070000",
         738 => x"13070000",
         739 => x"6ff01fef",
         740 => x"1307f000",
         741 => x"638ee700",
         742 => x"1307b000",
         743 => x"e382e7fc",
         744 => x"13880900",
         745 => x"13840400",
         746 => x"93060a00",
         747 => x"6ff09ffb",
         748 => x"37044000",
         749 => x"13080000",
         750 => x"93063000",
         751 => x"6ff09ffb",
         752 => x"93080900",
         753 => x"6ff01fe7",
         754 => x"93071000",
         755 => x"b387e740",
         756 => x"1307b001",
         757 => x"e348f7fa",
         758 => x"9388e809",
         759 => x"b357f400",
         760 => x"33141401",
         761 => x"33348000",
         762 => x"b3e78700",
         763 => x"13f77700",
         764 => x"630a0700",
         765 => x"13f7f700",
         766 => x"93064000",
         767 => x"6304d700",
         768 => x"93874700",
         769 => x"37070004",
         770 => x"33f7e700",
         771 => x"93d73700",
         772 => x"e30607e6",
         773 => x"93070000",
         774 => x"13071000",
         775 => x"6ff01fe6",
         776 => x"b7074000",
         777 => x"1307f00f",
         778 => x"13080000",
         779 => x"6ff01fe5",
         780 => x"93070000",
         781 => x"1307f00f",
         782 => x"6ff05fe4",
         783 => x"13060500",
         784 => x"13050000",
         785 => x"93f61500",
         786 => x"63840600",
         787 => x"3305c500",
         788 => x"93d51500",
         789 => x"13161600",
         790 => x"e39605fe",
         791 => x"67800000",
         792 => x"63400506",
         793 => x"63c60506",
         794 => x"13860500",
         795 => x"93050500",
         796 => x"1305f0ff",
         797 => x"630c0602",
         798 => x"93061000",
         799 => x"637ab600",
         800 => x"6358c000",
         801 => x"13161600",
         802 => x"93961600",
         803 => x"e36ab6fe",
         804 => x"13050000",
         805 => x"63e6c500",
         806 => x"b385c540",
         807 => x"3365d500",
         808 => x"93d61600",
         809 => x"13561600",
         810 => x"e39606fe",
         811 => x"67800000",
         812 => x"93820000",
         813 => x"eff05ffb",
         814 => x"13850500",
         815 => x"67800200",
         816 => x"3305a040",
         817 => x"6348b000",
         818 => x"b305b040",
         819 => x"6ff0dff9",
         820 => x"b305b040",
         821 => x"93820000",
         822 => x"eff01ff9",
         823 => x"3305a040",
         824 => x"67800200",
         825 => x"93820000",
         826 => x"63ca0500",
         827 => x"634c0500",
         828 => x"eff09ff7",
         829 => x"13850500",
         830 => x"67800200",
         831 => x"b305b040",
         832 => x"e35805fe",
         833 => x"3305a040",
         834 => x"eff01ff6",
         835 => x"3305b040",
         836 => x"67800200",
         837 => x"b7070100",
         838 => x"637af502",
         839 => x"93370510",
         840 => x"93c71700",
         841 => x"93973700",
         842 => x"37170000",
         843 => x"93060002",
         844 => x"b386f640",
         845 => x"3355f500",
         846 => x"930707f1",
         847 => x"b387a700",
         848 => x"03c50700",
         849 => x"3385a640",
         850 => x"67800000",
         851 => x"37070001",
         852 => x"93070001",
         853 => x"e36ae5fc",
         854 => x"93078001",
         855 => x"6ff0dffc",
         856 => x"b7170000",
         857 => x"83a70701",
         858 => x"130101fe",
         859 => x"37170000",
         860 => x"2326f100",
         861 => x"0325c100",
         862 => x"83254701",
         863 => x"232e1100",
         864 => x"eff04fb6",
         865 => x"2326a100",
         866 => x"b7170000",
         867 => x"0325c100",
         868 => x"83a58701",
         869 => x"eff04ffa",
         870 => x"2326a100",
         871 => x"b7170000",
         872 => x"0325c100",
         873 => x"83a5c701",
         874 => x"eff0dfb1",
         875 => x"8320c101",
         876 => x"2326a100",
         877 => x"13050000",
         878 => x"13010102",
         879 => x"67800000",
         880 => x"130101ff",
         881 => x"23248100",
         882 => x"23261100",
         883 => x"93070000",
         884 => x"13040500",
         885 => x"63880700",
         886 => x"93050000",
         887 => x"97000000",
         888 => x"e7000000",
         889 => x"b7170000",
         890 => x"03a50702",
         891 => x"83278502",
         892 => x"63840700",
         893 => x"e7800700",
         894 => x"13050400",
         895 => x"ef00000a",
         896 => x"130101ff",
         897 => x"23248100",
         898 => x"23229100",
         899 => x"37140000",
         900 => x"b7140000",
         901 => x"93874402",
         902 => x"13044402",
         903 => x"3304f440",
         904 => x"23202101",
         905 => x"23261100",
         906 => x"13542440",
         907 => x"93844402",
         908 => x"13090000",
         909 => x"63108904",
         910 => x"b7140000",
         911 => x"37140000",
         912 => x"93874402",
         913 => x"13044402",
         914 => x"3304f440",
         915 => x"13542440",
         916 => x"93844402",
         917 => x"13090000",
         918 => x"63188902",
         919 => x"8320c100",
         920 => x"03248100",
         921 => x"83244100",
         922 => x"03290100",
         923 => x"13010101",
         924 => x"67800000",
         925 => x"83a70400",
         926 => x"13091900",
         927 => x"93844400",
         928 => x"e7800700",
         929 => x"6ff01ffb",
         930 => x"83a70400",
         931 => x"13091900",
         932 => x"93844400",
         933 => x"e7800700",
         934 => x"6ff01ffc",
         935 => x"9308d005",
         936 => x"73000000",
         937 => x"63520502",
         938 => x"130101ff",
         939 => x"23248100",
         940 => x"13040500",
         941 => x"23261100",
         942 => x"33048040",
         943 => x"ef000001",
         944 => x"23208500",
         945 => x"6f000000",
         946 => x"6f000000",
         947 => x"03a50186",
         948 => x"67800000",
         949 => x"2c080000",
         950 => x"b8080000",
         951 => x"38080000",
         952 => x"b8080000",
         953 => x"a8080000",
         954 => x"b8080000",
         955 => x"38080000",
         956 => x"2c080000",
         957 => x"2c080000",
         958 => x"a8080000",
         959 => x"38080000",
         960 => x"08080000",
         961 => x"08080000",
         962 => x"08080000",
         963 => x"40080000",
         964 => x"00010202",
         965 => x"03030303",
         966 => x"04040404",
         967 => x"04040404",
         968 => x"05050505",
         969 => x"05050505",
         970 => x"05050505",
         971 => x"05050505",
         972 => x"06060606",
         973 => x"06060606",
         974 => x"06060606",
         975 => x"06060606",
         976 => x"06060606",
         977 => x"06060606",
         978 => x"06060606",
         979 => x"06060606",
         980 => x"07070707",
         981 => x"07070707",
         982 => x"07070707",
         983 => x"07070707",
         984 => x"07070707",
         985 => x"07070707",
         986 => x"07070707",
         987 => x"07070707",
         988 => x"07070707",
         989 => x"07070707",
         990 => x"07070707",
         991 => x"07070707",
         992 => x"07070707",
         993 => x"07070707",
         994 => x"07070707",
         995 => x"07070707",
         996 => x"08080808",
         997 => x"08080808",
         998 => x"08080808",
         999 => x"08080808",
        1000 => x"08080808",
        1001 => x"08080808",
        1002 => x"08080808",
        1003 => x"08080808",
        1004 => x"08080808",
        1005 => x"08080808",
        1006 => x"08080808",
        1007 => x"08080808",
        1008 => x"08080808",
        1009 => x"08080808",
        1010 => x"08080808",
        1011 => x"08080808",
        1012 => x"08080808",
        1013 => x"08080808",
        1014 => x"08080808",
        1015 => x"08080808",
        1016 => x"08080808",
        1017 => x"08080808",
        1018 => x"08080808",
        1019 => x"08080808",
        1020 => x"08080808",
        1021 => x"08080808",
        1022 => x"08080808",
        1023 => x"08080808",
        1024 => x"08080808",
        1025 => x"08080808",
        1026 => x"08080808",
        1027 => x"08080808",
        1028 => x"0000803f",
        1029 => x"00000040",
        1030 => x"000040c0",
        1031 => x"0000c8c1",
        1032 => x"00000020",
        1033 => x"00000000",
        1034 => x"00000000",
        1035 => x"00000000",
        1036 => x"00000000",
        1037 => x"00000000",
        1038 => x"00000000",
        1039 => x"00000000",
        1040 => x"00000000",
        1041 => x"00000000",
        1042 => x"00000000",
        1043 => x"00000000",
        1044 => x"00000000",
        1045 => x"00000000",
        1046 => x"00000000",
        1047 => x"00000000",
        1048 => x"00000000",
        1049 => x"00000000",
        1050 => x"00000000",
        1051 => x"00000000",
        1052 => x"00000000",
        1053 => x"00000000",
        1054 => x"00000000",
        1055 => x"00000000",
        1056 => x"00000000",
        1057 => x"00000020",
        others => (others => '-')
    );
end package processor_common_rom;
