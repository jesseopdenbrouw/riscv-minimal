-- srec2vhdl table generator
-- for input file string.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97",    1 => x"11",    2 => x"00",    3 => x"20", 
           4 => x"93",    5 => x"81",    6 => x"01",    7 => x"87", 
           8 => x"17",    9 => x"41",   10 => x"00",   11 => x"20", 
          12 => x"13",   13 => x"01",   14 => x"81",   15 => x"ff", 
          16 => x"33",   17 => x"04",   18 => x"01",   19 => x"00", 
          20 => x"b7",   21 => x"07",   22 => x"00",   23 => x"20", 
          24 => x"93",   25 => x"80",   26 => x"47",   27 => x"06", 
          28 => x"b7",   29 => x"07",   30 => x"00",   31 => x"20", 
          32 => x"93",   33 => x"84",   34 => x"47",   35 => x"06", 
          36 => x"13",   37 => x"09",   38 => x"40",   39 => x"25", 
          40 => x"6f",   41 => x"00",   42 => x"40",   43 => x"01", 
          44 => x"23",   45 => x"a0",   46 => x"00",   47 => x"00", 
          48 => x"93",   49 => x"87",   50 => x"00",   51 => x"00", 
          52 => x"93",   53 => x"80",   54 => x"47",   55 => x"00", 
          56 => x"83",   57 => x"a7",   58 => x"07",   59 => x"00", 
          60 => x"e3",   61 => x"e8",   62 => x"90",   63 => x"fe", 
          64 => x"b7",   65 => x"07",   66 => x"00",   67 => x"20", 
          68 => x"93",   69 => x"80",   70 => x"07",   71 => x"00", 
          72 => x"b7",   73 => x"07",   74 => x"00",   75 => x"20", 
          76 => x"93",   77 => x"84",   78 => x"07",   79 => x"06", 
          80 => x"6f",   81 => x"00",   82 => x"40",   83 => x"01", 
          84 => x"83",   85 => x"27",   86 => x"09",   87 => x"00", 
          88 => x"23",   89 => x"a0",   90 => x"f0",   91 => x"00", 
          92 => x"93",   93 => x"80",   94 => x"40",   95 => x"00", 
          96 => x"13",   97 => x"09",   98 => x"49",   99 => x"00", 
         100 => x"e3",  101 => x"e8",  102 => x"90",  103 => x"fe", 
         104 => x"ef",  105 => x"00",  106 => x"00",  107 => x"0d", 
         108 => x"ef",  109 => x"00",  110 => x"c0",  111 => x"00", 
         112 => x"13",  113 => x"05",  114 => x"00",  115 => x"00", 
         116 => x"ef",  117 => x"00",  118 => x"80",  119 => x"08", 
         120 => x"13",  121 => x"01",  122 => x"01",  123 => x"f7", 
         124 => x"23",  125 => x"26",  126 => x"11",  127 => x"08", 
         128 => x"23",  129 => x"24",  130 => x"81",  131 => x"08", 
         132 => x"13",  133 => x"04",  134 => x"01",  135 => x"09", 
         136 => x"93",  137 => x"07",  138 => x"80",  139 => x"23", 
         140 => x"03",  141 => x"a5",  142 => x"07",  143 => x"00", 
         144 => x"83",  145 => x"a5",  146 => x"47",  147 => x"00", 
         148 => x"03",  149 => x"a6",  150 => x"87",  151 => x"00", 
         152 => x"83",  153 => x"a6",  154 => x"c7",  155 => x"00", 
         156 => x"03",  157 => x"a7",  158 => x"07",  159 => x"01", 
         160 => x"83",  161 => x"a7",  162 => x"47",  163 => x"01", 
         164 => x"23",  165 => x"2c",  166 => x"a4",  167 => x"fc", 
         168 => x"23",  169 => x"2e",  170 => x"b4",  171 => x"fc", 
         172 => x"23",  173 => x"20",  174 => x"c4",  175 => x"fe", 
         176 => x"23",  177 => x"22",  178 => x"d4",  179 => x"fe", 
         180 => x"23",  181 => x"24",  182 => x"e4",  183 => x"fe", 
         184 => x"23",  185 => x"26",  186 => x"f4",  187 => x"fe", 
         188 => x"93",  189 => x"07",  190 => x"84",  191 => x"fd", 
         192 => x"13",  193 => x"85",  194 => x"07",  195 => x"00", 
         196 => x"ef",  197 => x"00",  198 => x"c0",  199 => x"11", 
         200 => x"93",  201 => x"07",  202 => x"05",  203 => x"00", 
         204 => x"23",  205 => x"28",  206 => x"f4",  207 => x"f6", 
         208 => x"13",  209 => x"07",  210 => x"84",  211 => x"fd", 
         212 => x"93",  213 => x"07",  214 => x"44",  215 => x"f7", 
         216 => x"93",  217 => x"05",  218 => x"07",  219 => x"00", 
         220 => x"13",  221 => x"85",  222 => x"07",  223 => x"00", 
         224 => x"ef",  225 => x"00",  226 => x"40",  227 => x"0e", 
         228 => x"83",  229 => x"27",  230 => x"04",  231 => x"f7", 
         232 => x"13",  233 => x"85",  234 => x"07",  235 => x"00", 
         236 => x"83",  237 => x"20",  238 => x"c1",  239 => x"08", 
         240 => x"03",  241 => x"24",  242 => x"81",  243 => x"08", 
         244 => x"13",  245 => x"01",  246 => x"01",  247 => x"09", 
         248 => x"67",  249 => x"80",  250 => x"00",  251 => x"00", 
         252 => x"13",  253 => x"01",  254 => x"01",  255 => x"ff", 
         256 => x"23",  257 => x"24",  258 => x"81",  259 => x"00", 
         260 => x"23",  261 => x"26",  262 => x"11",  263 => x"00", 
         264 => x"93",  265 => x"07",  266 => x"00",  267 => x"00", 
         268 => x"13",  269 => x"04",  270 => x"05",  271 => x"00", 
         272 => x"63",  273 => x"88",  274 => x"07",  275 => x"00", 
         276 => x"93",  277 => x"05",  278 => x"00",  279 => x"00", 
         280 => x"97",  281 => x"00",  282 => x"00",  283 => x"00", 
         284 => x"e7",  285 => x"00",  286 => x"00",  287 => x"00", 
         288 => x"03",  289 => x"25",  290 => x"00",  291 => x"25", 
         292 => x"83",  293 => x"27",  294 => x"85",  295 => x"02", 
         296 => x"63",  297 => x"84",  298 => x"07",  299 => x"00", 
         300 => x"e7",  301 => x"80",  302 => x"07",  303 => x"00", 
         304 => x"13",  305 => x"05",  306 => x"04",  307 => x"00", 
         308 => x"ef",  309 => x"00",  310 => x"80",  311 => x"0c", 
         312 => x"13",  313 => x"01",  314 => x"01",  315 => x"ff", 
         316 => x"23",  317 => x"24",  318 => x"81",  319 => x"00", 
         320 => x"23",  321 => x"22",  322 => x"91",  323 => x"00", 
         324 => x"93",  325 => x"07",  326 => x"40",  327 => x"25", 
         328 => x"13",  329 => x"04",  330 => x"40",  331 => x"25", 
         332 => x"33",  333 => x"04",  334 => x"f4",  335 => x"40", 
         336 => x"23",  337 => x"20",  338 => x"21",  339 => x"01", 
         340 => x"23",  341 => x"26",  342 => x"11",  343 => x"00", 
         344 => x"13",  345 => x"54",  346 => x"24",  347 => x"40", 
         348 => x"93",  349 => x"04",  350 => x"40",  351 => x"25", 
         352 => x"13",  353 => x"09",  354 => x"00",  355 => x"00", 
         356 => x"63",  357 => x"1c",  358 => x"89",  359 => x"02", 
         360 => x"93",  361 => x"07",  362 => x"40",  363 => x"25", 
         364 => x"13",  365 => x"04",  366 => x"40",  367 => x"25", 
         368 => x"33",  369 => x"04",  370 => x"f4",  371 => x"40", 
         372 => x"13",  373 => x"54",  374 => x"24",  375 => x"40", 
         376 => x"93",  377 => x"04",  378 => x"40",  379 => x"25", 
         380 => x"13",  381 => x"09",  382 => x"00",  383 => x"00", 
         384 => x"63",  385 => x"18",  386 => x"89",  387 => x"02", 
         388 => x"83",  389 => x"20",  390 => x"c1",  391 => x"00", 
         392 => x"03",  393 => x"24",  394 => x"81",  395 => x"00", 
         396 => x"83",  397 => x"24",  398 => x"41",  399 => x"00", 
         400 => x"03",  401 => x"29",  402 => x"01",  403 => x"00", 
         404 => x"13",  405 => x"01",  406 => x"01",  407 => x"01", 
         408 => x"67",  409 => x"80",  410 => x"00",  411 => x"00", 
         412 => x"83",  413 => x"a7",  414 => x"04",  415 => x"00", 
         416 => x"13",  417 => x"09",  418 => x"19",  419 => x"00", 
         420 => x"93",  421 => x"84",  422 => x"44",  423 => x"00", 
         424 => x"e7",  425 => x"80",  426 => x"07",  427 => x"00", 
         428 => x"6f",  429 => x"f0",  430 => x"9f",  431 => x"fb", 
         432 => x"83",  433 => x"a7",  434 => x"04",  435 => x"00", 
         436 => x"13",  437 => x"09",  438 => x"19",  439 => x"00", 
         440 => x"93",  441 => x"84",  442 => x"44",  443 => x"00", 
         444 => x"e7",  445 => x"80",  446 => x"07",  447 => x"00", 
         448 => x"6f",  449 => x"f0",  450 => x"1f",  451 => x"fc", 
         452 => x"93",  453 => x"07",  454 => x"05",  455 => x"00", 
         456 => x"03",  457 => x"c7",  458 => x"05",  459 => x"00", 
         460 => x"93",  461 => x"87",  462 => x"17",  463 => x"00", 
         464 => x"93",  465 => x"85",  466 => x"15",  467 => x"00", 
         468 => x"a3",  469 => x"8f",  470 => x"e7",  471 => x"fe", 
         472 => x"e3",  473 => x"18",  474 => x"07",  475 => x"fe", 
         476 => x"67",  477 => x"80",  478 => x"00",  479 => x"00", 
         480 => x"93",  481 => x"07",  482 => x"05",  483 => x"00", 
         484 => x"03",  485 => x"c7",  486 => x"07",  487 => x"00", 
         488 => x"93",  489 => x"87",  490 => x"17",  491 => x"00", 
         492 => x"e3",  493 => x"1c",  494 => x"07",  495 => x"fe", 
         496 => x"33",  497 => x"85",  498 => x"a7",  499 => x"40", 
         500 => x"13",  501 => x"05",  502 => x"f5",  503 => x"ff", 
         504 => x"67",  505 => x"80",  506 => x"00",  507 => x"00", 
         508 => x"93",  509 => x"08",  510 => x"d0",  511 => x"05", 
         512 => x"73",  513 => x"00",  514 => x"00",  515 => x"00", 
         516 => x"63",  517 => x"52",  518 => x"05",  519 => x"02", 
         520 => x"13",  521 => x"01",  522 => x"01",  523 => x"ff", 
         524 => x"23",  525 => x"24",  526 => x"81",  527 => x"00", 
         528 => x"13",  529 => x"04",  530 => x"05",  531 => x"00", 
         532 => x"23",  533 => x"26",  534 => x"11",  535 => x"00", 
         536 => x"33",  537 => x"04",  538 => x"80",  539 => x"40", 
         540 => x"ef",  541 => x"00",  542 => x"00",  543 => x"01", 
         544 => x"23",  545 => x"20",  546 => x"85",  547 => x"00", 
         548 => x"6f",  549 => x"00",  550 => x"00",  551 => x"00", 
         552 => x"6f",  553 => x"00",  554 => x"00",  555 => x"00", 
         556 => x"b7",  557 => x"07",  558 => x"00",  559 => x"20", 
         560 => x"03",  561 => x"a5",  562 => x"07",  563 => x"06", 
         564 => x"67",  565 => x"80",  566 => x"00",  567 => x"00", 
         568 => x"48",  569 => x"65",  570 => x"6c",  571 => x"6c", 
         572 => x"6f",  573 => x"20",  574 => x"64",  575 => x"69", 
         576 => x"74",  577 => x"20",  578 => x"69",  579 => x"73", 
         580 => x"20",  581 => x"65",  582 => x"65",  583 => x"6e", 
         584 => x"20",  585 => x"73",  586 => x"74",  587 => x"72", 
         588 => x"69",  589 => x"6e",  590 => x"67",  591 => x"00", 
         592 => x"00",  593 => x"00",  594 => x"00",  595 => x"20", 
         596 => x"00",  597 => x"00",  598 => x"00",  599 => x"00", 
         600 => x"00",  601 => x"00",  602 => x"00",  603 => x"00", 
         604 => x"00",  605 => x"00",  606 => x"00",  607 => x"00", 
         608 => x"00",  609 => x"00",  610 => x"00",  611 => x"00", 
         612 => x"00",  613 => x"00",  614 => x"00",  615 => x"00", 
         616 => x"00",  617 => x"00",  618 => x"00",  619 => x"00", 
         620 => x"00",  621 => x"00",  622 => x"00",  623 => x"00", 
         624 => x"00",  625 => x"00",  626 => x"00",  627 => x"00", 
         628 => x"00",  629 => x"00",  630 => x"00",  631 => x"00", 
         632 => x"00",  633 => x"00",  634 => x"00",  635 => x"00", 
         636 => x"00",  637 => x"00",  638 => x"00",  639 => x"00", 
         640 => x"00",  641 => x"00",  642 => x"00",  643 => x"00", 
         644 => x"00",  645 => x"00",  646 => x"00",  647 => x"00", 
         648 => x"00",  649 => x"00",  650 => x"00",  651 => x"00", 
         652 => x"00",  653 => x"00",  654 => x"00",  655 => x"00", 
         656 => x"00",  657 => x"00",  658 => x"00",  659 => x"00", 
         660 => x"00",  661 => x"00",  662 => x"00",  663 => x"00", 
         664 => x"00",  665 => x"00",  666 => x"00",  667 => x"00", 
         668 => x"00",  669 => x"00",  670 => x"00",  671 => x"00", 
         672 => x"00",  673 => x"00",  674 => x"00",  675 => x"00", 
         676 => x"00",  677 => x"00",  678 => x"00",  679 => x"00", 
         680 => x"00",  681 => x"00",  682 => x"00",  683 => x"00", 
         684 => x"00",  685 => x"00",  686 => x"00",  687 => x"00", 
         688 => x"00",  689 => x"00",  690 => x"00",  691 => x"00", 
         692 => x"00",  693 => x"00",  694 => x"00",  695 => x"20", 
        others => (others => '-')
    );
end package processor_common_rom;
