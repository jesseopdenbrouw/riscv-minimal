-- srec2vhdl table generator
-- for input file malloc.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"93804186",
           5 => x"93844187",
           6 => x"b7170000",
           7 => x"13894793",
           8 => x"6f004001",
           9 => x"23a00000",
          10 => x"93870000",
          11 => x"93804700",
          12 => x"83a70700",
          13 => x"e3e890fe",
          14 => x"b7070020",
          15 => x"93800700",
          16 => x"93844186",
          17 => x"6f004001",
          18 => x"83270900",
          19 => x"23a0f000",
          20 => x"93804000",
          21 => x"13094900",
          22 => x"e3e890fe",
          23 => x"ef00002b",
          24 => x"ef00c000",
          25 => x"13050000",
          26 => x"ef004026",
          27 => x"130101fd",
          28 => x"23261102",
          29 => x"23248102",
          30 => x"13040103",
          31 => x"13054006",
          32 => x"ef008032",
          33 => x"93070500",
          34 => x"232ef4fc",
          35 => x"232604fe",
          36 => x"6f004002",
          37 => x"8327c4fe",
          38 => x"0327c4fd",
          39 => x"b307f700",
          40 => x"13071004",
          41 => x"2380e700",
          42 => x"8327c4fe",
          43 => x"93871700",
          44 => x"2326f4fe",
          45 => x"0327c4fe",
          46 => x"93073006",
          47 => x"e3dce7fc",
          48 => x"0325c4fd",
          49 => x"ef00002f",
          50 => x"13052003",
          51 => x"ef00c02d",
          52 => x"93070500",
          53 => x"232ef4fc",
          54 => x"232404fe",
          55 => x"6f000003",
          56 => x"832784fe",
          57 => x"13f7f70f",
          58 => x"832784fe",
          59 => x"8326c4fd",
          60 => x"b387f600",
          61 => x"13071704",
          62 => x"1377f70f",
          63 => x"2380e700",
          64 => x"832784fe",
          65 => x"93871700",
          66 => x"2324f4fe",
          67 => x"032784fe",
          68 => x"93071003",
          69 => x"e3d6e7fc",
          70 => x"0325c4fd",
          71 => x"ef008029",
          72 => x"13054006",
          73 => x"ef004028",
          74 => x"93070500",
          75 => x"232cf4fc",
          76 => x"232204fe",
          77 => x"6f008002",
          78 => x"832744fe",
          79 => x"93972700",
          80 => x"032784fd",
          81 => x"b307f700",
          82 => x"1307f0ff",
          83 => x"23a0e700",
          84 => x"832744fe",
          85 => x"93871700",
          86 => x"2322f4fe",
          87 => x"032744fe",
          88 => x"93078001",
          89 => x"e3dae7fc",
          90 => x"032584fd",
          91 => x"ef008024",
          92 => x"93054000",
          93 => x"13059001",
          94 => x"ef00c013",
          95 => x"93070500",
          96 => x"232af4fc",
          97 => x"232004fe",
          98 => x"6f00c002",
          99 => x"832704fe",
         100 => x"93972700",
         101 => x"032744fd",
         102 => x"b307f700",
         103 => x"37171111",
         104 => x"13071711",
         105 => x"23a0e700",
         106 => x"832704fe",
         107 => x"93871700",
         108 => x"2320f4fe",
         109 => x"032704fe",
         110 => x"93078001",
         111 => x"e3d8e7fc",
         112 => x"93070000",
         113 => x"13850700",
         114 => x"8320c102",
         115 => x"03248102",
         116 => x"13010103",
         117 => x"67800000",
         118 => x"130101fd",
         119 => x"23261102",
         120 => x"23248102",
         121 => x"13040103",
         122 => x"232ea4fc",
         123 => x"b7870020",
         124 => x"13870700",
         125 => x"93070040",
         126 => x"b307f740",
         127 => x"2326f4fe",
         128 => x"8327c4fe",
         129 => x"2324f4fe",
         130 => x"83a70187",
         131 => x"63960700",
         132 => x"13878187",
         133 => x"23a8e186",
         134 => x"03a70187",
         135 => x"8327c4fd",
         136 => x"b307f700",
         137 => x"032784fe",
         138 => x"637ef700",
         139 => x"ef008009",
         140 => x"13070500",
         141 => x"9307c000",
         142 => x"2320f700",
         143 => x"9307f0ff",
         144 => x"6f000002",
         145 => x"83a70187",
         146 => x"2322f4fe",
         147 => x"03a70187",
         148 => x"8327c4fd",
         149 => x"3307f700",
         150 => x"23a8e186",
         151 => x"832744fe",
         152 => x"13850700",
         153 => x"8320c102",
         154 => x"03248102",
         155 => x"13010103",
         156 => x"67800000",
         157 => x"13030500",
         158 => x"630a0600",
         159 => x"2300b300",
         160 => x"1306f6ff",
         161 => x"13031300",
         162 => x"e31a06fe",
         163 => x"67800000",
         164 => x"13060500",
         165 => x"13050000",
         166 => x"93f61500",
         167 => x"63840600",
         168 => x"3305c500",
         169 => x"93d51500",
         170 => x"13161600",
         171 => x"e39605fe",
         172 => x"67800000",
         173 => x"13860500",
         174 => x"93050500",
         175 => x"03a50186",
         176 => x"6f000010",
         177 => x"03a50186",
         178 => x"67800000",
         179 => x"130101ff",
         180 => x"23248100",
         181 => x"23261100",
         182 => x"93070000",
         183 => x"13040500",
         184 => x"63880700",
         185 => x"93050000",
         186 => x"97000000",
         187 => x"e7000000",
         188 => x"b7170000",
         189 => x"03a50793",
         190 => x"83278502",
         191 => x"63840700",
         192 => x"e7800700",
         193 => x"13050400",
         194 => x"ef00805f",
         195 => x"130101ff",
         196 => x"23248100",
         197 => x"23229100",
         198 => x"37140000",
         199 => x"b7140000",
         200 => x"93874493",
         201 => x"13044493",
         202 => x"3304f440",
         203 => x"23202101",
         204 => x"23261100",
         205 => x"13542440",
         206 => x"93844493",
         207 => x"13090000",
         208 => x"63108904",
         209 => x"b7140000",
         210 => x"37140000",
         211 => x"93874493",
         212 => x"13044493",
         213 => x"3304f440",
         214 => x"13542440",
         215 => x"93844493",
         216 => x"13090000",
         217 => x"63188902",
         218 => x"8320c100",
         219 => x"03248100",
         220 => x"83244100",
         221 => x"03290100",
         222 => x"13010101",
         223 => x"67800000",
         224 => x"83a70400",
         225 => x"13091900",
         226 => x"93844400",
         227 => x"e7800700",
         228 => x"6ff01ffb",
         229 => x"83a70400",
         230 => x"13091900",
         231 => x"93844400",
         232 => x"e7800700",
         233 => x"6ff01ffc",
         234 => x"93050500",
         235 => x"03a50186",
         236 => x"6f008020",
         237 => x"93050500",
         238 => x"03a50186",
         239 => x"6f004010",
         240 => x"130101fd",
         241 => x"23229102",
         242 => x"23202103",
         243 => x"23261102",
         244 => x"23248102",
         245 => x"232e3101",
         246 => x"13d90501",
         247 => x"93040500",
         248 => x"93560601",
         249 => x"13850500",
         250 => x"6310090a",
         251 => x"63920604",
         252 => x"93150601",
         253 => x"13150501",
         254 => x"93d50501",
         255 => x"13550501",
         256 => x"eff01fe9",
         257 => x"13060500",
         258 => x"93050600",
         259 => x"13850400",
         260 => x"2326c100",
         261 => x"ef00401a",
         262 => x"13040500",
         263 => x"63020508",
         264 => x"0326c100",
         265 => x"93050000",
         266 => x"eff0dfe4",
         267 => x"6f004007",
         268 => x"13890600",
         269 => x"93890500",
         270 => x"93150601",
         271 => x"13150501",
         272 => x"93d50501",
         273 => x"13550501",
         274 => x"eff09fe4",
         275 => x"13040500",
         276 => x"93150901",
         277 => x"13950901",
         278 => x"93d50501",
         279 => x"13550501",
         280 => x"eff01fe3",
         281 => x"93570401",
         282 => x"3306f500",
         283 => x"93570601",
         284 => x"63920702",
         285 => x"13140401",
         286 => x"13160601",
         287 => x"13540401",
         288 => x"33668600",
         289 => x"6ff05ff8",
         290 => x"63960600",
         291 => x"93090600",
         292 => x"6ff09ffa",
         293 => x"9307c000",
         294 => x"23a0f400",
         295 => x"13040000",
         296 => x"8320c102",
         297 => x"13050400",
         298 => x"03248102",
         299 => x"83244102",
         300 => x"03290102",
         301 => x"8329c101",
         302 => x"13010103",
         303 => x"67800000",
         304 => x"638a050e",
         305 => x"83a7c5ff",
         306 => x"130101fe",
         307 => x"232c8100",
         308 => x"232e1100",
         309 => x"1384c5ff",
         310 => x"63d40700",
         311 => x"3304f400",
         312 => x"2326a100",
         313 => x"ef00c026",
         314 => x"83a74186",
         315 => x"0325c100",
         316 => x"639e0700",
         317 => x"23220400",
         318 => x"23a28186",
         319 => x"03248101",
         320 => x"8320c101",
         321 => x"13010102",
         322 => x"6f00c024",
         323 => x"6374f402",
         324 => x"03260400",
         325 => x"b306c400",
         326 => x"639ad700",
         327 => x"83a60700",
         328 => x"83a74700",
         329 => x"b386c600",
         330 => x"2320d400",
         331 => x"2322f400",
         332 => x"6ff09ffc",
         333 => x"13870700",
         334 => x"83a74700",
         335 => x"63840700",
         336 => x"e37af4fe",
         337 => x"83260700",
         338 => x"3306d700",
         339 => x"63188602",
         340 => x"03260400",
         341 => x"b386c600",
         342 => x"2320d700",
         343 => x"3306d700",
         344 => x"e39ec7f8",
         345 => x"03a60700",
         346 => x"83a74700",
         347 => x"b306d600",
         348 => x"2320d700",
         349 => x"2322f700",
         350 => x"6ff05ff8",
         351 => x"6378c400",
         352 => x"9307c000",
         353 => x"2320f500",
         354 => x"6ff05ff7",
         355 => x"03260400",
         356 => x"b306c400",
         357 => x"639ad700",
         358 => x"83a60700",
         359 => x"83a74700",
         360 => x"b386c600",
         361 => x"2320d400",
         362 => x"2322f400",
         363 => x"23228700",
         364 => x"6ff0dff4",
         365 => x"67800000",
         366 => x"130101fe",
         367 => x"232a9100",
         368 => x"93843500",
         369 => x"93f4c4ff",
         370 => x"23282101",
         371 => x"232e1100",
         372 => x"232c8100",
         373 => x"23263101",
         374 => x"93848400",
         375 => x"9307c000",
         376 => x"13090500",
         377 => x"63f4f406",
         378 => x"9304c000",
         379 => x"63e2b406",
         380 => x"13050900",
         381 => x"ef00c015",
         382 => x"03a74186",
         383 => x"93864186",
         384 => x"13040700",
         385 => x"631a0406",
         386 => x"13848186",
         387 => x"83270400",
         388 => x"639a0700",
         389 => x"93050000",
         390 => x"13050900",
         391 => x"ef00c00e",
         392 => x"2320a400",
         393 => x"93850400",
         394 => x"13050900",
         395 => x"ef00c00d",
         396 => x"9309f0ff",
         397 => x"631a350b",
         398 => x"9307c000",
         399 => x"2320f900",
         400 => x"13050900",
         401 => x"ef000011",
         402 => x"6f000001",
         403 => x"e3d004fa",
         404 => x"9307c000",
         405 => x"2320f900",
         406 => x"13050000",
         407 => x"8320c101",
         408 => x"03248101",
         409 => x"83244101",
         410 => x"03290101",
         411 => x"8329c100",
         412 => x"13010102",
         413 => x"67800000",
         414 => x"83270400",
         415 => x"b3879740",
         416 => x"63ce0704",
         417 => x"1306b000",
         418 => x"637af600",
         419 => x"2320f400",
         420 => x"3304f400",
         421 => x"23209400",
         422 => x"6f000001",
         423 => x"83274400",
         424 => x"631a8702",
         425 => x"23a0f600",
         426 => x"13050900",
         427 => x"ef00800a",
         428 => x"1305b400",
         429 => x"93074400",
         430 => x"137585ff",
         431 => x"3307f540",
         432 => x"e30ef5f8",
         433 => x"3304e400",
         434 => x"b387a740",
         435 => x"2320f400",
         436 => x"6ff0dff8",
         437 => x"2322f700",
         438 => x"6ff01ffd",
         439 => x"13070400",
         440 => x"03244400",
         441 => x"6ff01ff2",
         442 => x"13043500",
         443 => x"1374c4ff",
         444 => x"e30285fa",
         445 => x"b305a440",
         446 => x"13050900",
         447 => x"ef00c000",
         448 => x"e31a35f9",
         449 => x"6ff05ff3",
         450 => x"130101ff",
         451 => x"23248100",
         452 => x"23229100",
         453 => x"13040500",
         454 => x"13850500",
         455 => x"23261100",
         456 => x"23a60186",
         457 => x"eff05fab",
         458 => x"9307f0ff",
         459 => x"6318f500",
         460 => x"83a7c186",
         461 => x"63840700",
         462 => x"2320f400",
         463 => x"8320c100",
         464 => x"03248100",
         465 => x"83244100",
         466 => x"13010101",
         467 => x"67800000",
         468 => x"67800000",
         469 => x"67800000",
         470 => x"130101ff",
         471 => x"23248100",
         472 => x"13840500",
         473 => x"83a50500",
         474 => x"23229100",
         475 => x"23261100",
         476 => x"93040500",
         477 => x"63840500",
         478 => x"eff01ffe",
         479 => x"93050400",
         480 => x"03248100",
         481 => x"8320c100",
         482 => x"13850400",
         483 => x"83244100",
         484 => x"13010101",
         485 => x"6ff0dfd2",
         486 => x"83a70186",
         487 => x"6380a716",
         488 => x"83274502",
         489 => x"130101fe",
         490 => x"232c8100",
         491 => x"232e1100",
         492 => x"232a9100",
         493 => x"23282101",
         494 => x"23263101",
         495 => x"13040500",
         496 => x"63840702",
         497 => x"83a7c700",
         498 => x"93040000",
         499 => x"13090008",
         500 => x"6392070e",
         501 => x"83274402",
         502 => x"83a50700",
         503 => x"63860500",
         504 => x"13050400",
         505 => x"eff0dfcd",
         506 => x"83254401",
         507 => x"63860500",
         508 => x"13050400",
         509 => x"eff0dfcc",
         510 => x"83254402",
         511 => x"63860500",
         512 => x"13050400",
         513 => x"eff0dfcb",
         514 => x"83258403",
         515 => x"63860500",
         516 => x"13050400",
         517 => x"eff0dfca",
         518 => x"8325c403",
         519 => x"63860500",
         520 => x"13050400",
         521 => x"eff0dfc9",
         522 => x"83250404",
         523 => x"63860500",
         524 => x"13050400",
         525 => x"eff0dfc8",
         526 => x"8325c405",
         527 => x"63860500",
         528 => x"13050400",
         529 => x"eff0dfc7",
         530 => x"83258405",
         531 => x"63860500",
         532 => x"13050400",
         533 => x"eff0dfc6",
         534 => x"83254403",
         535 => x"63860500",
         536 => x"13050400",
         537 => x"eff0dfc5",
         538 => x"83278401",
         539 => x"638a0706",
         540 => x"83278402",
         541 => x"13050400",
         542 => x"e7800700",
         543 => x"83258404",
         544 => x"63800506",
         545 => x"13050400",
         546 => x"03248101",
         547 => x"8320c101",
         548 => x"83244101",
         549 => x"03290101",
         550 => x"8329c100",
         551 => x"13010102",
         552 => x"6ff09feb",
         553 => x"b3859500",
         554 => x"83a50500",
         555 => x"63900502",
         556 => x"93844400",
         557 => x"83274402",
         558 => x"83a5c700",
         559 => x"e39424ff",
         560 => x"13050400",
         561 => x"eff0dfbf",
         562 => x"6ff0dff0",
         563 => x"83a90500",
         564 => x"13050400",
         565 => x"eff0dfbe",
         566 => x"93850900",
         567 => x"6ff01ffd",
         568 => x"8320c101",
         569 => x"03248101",
         570 => x"83244101",
         571 => x"03290101",
         572 => x"8329c100",
         573 => x"13010102",
         574 => x"67800000",
         575 => x"67800000",
         576 => x"9308d005",
         577 => x"73000000",
         578 => x"63520502",
         579 => x"130101ff",
         580 => x"23248100",
         581 => x"13040500",
         582 => x"23261100",
         583 => x"33048040",
         584 => x"eff05f9a",
         585 => x"23208500",
         586 => x"6f000000",
         587 => x"6f000000",
         588 => x"00000020",
         589 => x"00000000",
         590 => x"00000000",
         591 => x"00000000",
         592 => x"00000000",
         593 => x"00000000",
         594 => x"00000000",
         595 => x"00000000",
         596 => x"00000000",
         597 => x"00000000",
         598 => x"00000000",
         599 => x"00000000",
         600 => x"00000000",
         601 => x"00000000",
         602 => x"00000000",
         603 => x"00000000",
         604 => x"00000000",
         605 => x"00000000",
         606 => x"00000000",
         607 => x"00000000",
         608 => x"00000000",
         609 => x"00000000",
         610 => x"00000000",
         611 => x"00000000",
         612 => x"00000000",
         613 => x"00000020",
        others => (others => '0')
    );
end package processor_common_rom;
