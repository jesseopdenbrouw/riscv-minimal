-- srec2vhdl table generator
-- for input file main.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"93828206",
           6 => x"73905230",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef109008",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"9385c537",
          21 => x"13050500",
          22 => x"ef101004",
          23 => x"ef10902a",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10500a",
          29 => x"ef101025",
          30 => x"6f000000",
          31 => x"b70700f0",
          32 => x"1307101b",
          33 => x"23a2e702",
          34 => x"13070004",
          35 => x"23a4e702",
          36 => x"67800000",
          37 => x"1375f50f",
          38 => x"b70700f0",
          39 => x"23a0a702",
          40 => x"370700f0",
          41 => x"8327c702",
          42 => x"93f70701",
          43 => x"e38c07fe",
          44 => x"67800000",
          45 => x"63060502",
          46 => x"83470500",
          47 => x"63820702",
          48 => x"370700f0",
          49 => x"13051500",
          50 => x"2320f702",
          51 => x"8327c702",
          52 => x"93f70701",
          53 => x"e38c07fe",
          54 => x"83470500",
          55 => x"e39407fe",
          56 => x"67800000",
          57 => x"370700f0",
          58 => x"8327c702",
          59 => x"93f74700",
          60 => x"e38c07fe",
          61 => x"03250702",
          62 => x"1375f50f",
          63 => x"67800000",
          64 => x"130101ff",
          65 => x"373e0000",
          66 => x"370700f0",
          67 => x"930e0500",
          68 => x"138ff5ff",
          69 => x"23268100",
          70 => x"13050000",
          71 => x"130e8efb",
          72 => x"13070702",
          73 => x"13035001",
          74 => x"93027000",
          75 => x"930fe005",
          76 => x"9305f007",
          77 => x"93082000",
          78 => x"13082001",
          79 => x"b7330000",
          80 => x"1306f007",
          81 => x"8327c700",
          82 => x"93f74700",
          83 => x"e38c07fe",
          84 => x"03240700",
          85 => x"9376f40f",
          86 => x"636ed302",
          87 => x"63fed802",
          88 => x"9387d6ff",
          89 => x"636af802",
          90 => x"93972700",
          91 => x"b307fe00",
          92 => x"83a70700",
          93 => x"67800700",
          94 => x"1305f5ff",
          95 => x"6308050c",
          96 => x"2320c700",
          97 => x"8327c700",
          98 => x"93f70701",
          99 => x"e38c07fe",
         100 => x"6ff09ffe",
         101 => x"638cb606",
         102 => x"635ae50d",
         103 => x"1374f40f",
         104 => x"930704fe",
         105 => x"93f7f70f",
         106 => x"e3eefff8",
         107 => x"b387ae00",
         108 => x"23808700",
         109 => x"13051500",
         110 => x"2320d700",
         111 => x"8327c700",
         112 => x"93f70701",
         113 => x"e38c07fe",
         114 => x"6ff0dff7",
         115 => x"b38eae00",
         116 => x"b7360000",
         117 => x"23800e00",
         118 => x"9307d000",
         119 => x"93864620",
         120 => x"370700f0",
         121 => x"93861600",
         122 => x"2320f702",
         123 => x"8327c702",
         124 => x"93f70701",
         125 => x"e38c07fe",
         126 => x"83c70600",
         127 => x"e39407fe",
         128 => x"0324c100",
         129 => x"13010101",
         130 => x"67800000",
         131 => x"63040504",
         132 => x"2320b700",
         133 => x"8327c700",
         134 => x"93f70701",
         135 => x"e38c07fe",
         136 => x"1305f5ff",
         137 => x"6ff01ff2",
         138 => x"9307c003",
         139 => x"9386432c",
         140 => x"93861600",
         141 => x"2320f700",
         142 => x"8327c700",
         143 => x"93f70701",
         144 => x"e38c07fe",
         145 => x"83c70600",
         146 => x"e39407fe",
         147 => x"13050000",
         148 => x"6ff05fef",
         149 => x"23205700",
         150 => x"8327c700",
         151 => x"93f70701",
         152 => x"e38c07fe",
         153 => x"13050000",
         154 => x"6ff0dfed",
         155 => x"23205700",
         156 => x"8327c700",
         157 => x"93f70701",
         158 => x"e38c07fe",
         159 => x"6ff09fec",
         160 => x"1375f50f",
         161 => x"b70700f0",
         162 => x"23a0a702",
         163 => x"370700f0",
         164 => x"8327c702",
         165 => x"93f70701",
         166 => x"e38c07fe",
         167 => x"13051000",
         168 => x"67800000",
         169 => x"370700f0",
         170 => x"8327c702",
         171 => x"93f74700",
         172 => x"e38c07fe",
         173 => x"03250702",
         174 => x"1375f50f",
         175 => x"67800000",
         176 => x"13050000",
         177 => x"67800000",
         178 => x"13050000",
         179 => x"67800000",
         180 => x"6f000008",
         181 => x"6f004043",
         182 => x"6f000043",
         183 => x"6f00c042",
         184 => x"6f008042",
         185 => x"6f004042",
         186 => x"6f000042",
         187 => x"6f000042",
         188 => x"6f008041",
         189 => x"6f004041",
         190 => x"6f000041",
         191 => x"6f00c040",
         192 => x"6f008040",
         193 => x"6f004040",
         194 => x"6f000040",
         195 => x"6f00c03f",
         196 => x"6f00803f",
         197 => x"6f00403b",
         198 => x"6f008046",
         199 => x"6f00c03e",
         200 => x"6f00803e",
         201 => x"6f00403e",
         202 => x"6f00003e",
         203 => x"6f00c03d",
         204 => x"6f00803d",
         205 => x"6f00403d",
         206 => x"6f00003d",
         207 => x"6f00c03c",
         208 => x"6f00803c",
         209 => x"6f00403c",
         210 => x"6f00003c",
         211 => x"6f00c03b",
         212 => x"130101f8",
         213 => x"23221100",
         214 => x"23242100",
         215 => x"23263100",
         216 => x"23284100",
         217 => x"232a5100",
         218 => x"232c6100",
         219 => x"232e7100",
         220 => x"23208102",
         221 => x"23229102",
         222 => x"2324a102",
         223 => x"2326b102",
         224 => x"2328c102",
         225 => x"232ad102",
         226 => x"232ce102",
         227 => x"232ef102",
         228 => x"23200105",
         229 => x"23221105",
         230 => x"23242105",
         231 => x"23263105",
         232 => x"23284105",
         233 => x"232a5105",
         234 => x"232c6105",
         235 => x"232e7105",
         236 => x"23208107",
         237 => x"23229107",
         238 => x"2324a107",
         239 => x"2326b107",
         240 => x"2328c107",
         241 => x"232ad107",
         242 => x"232ce107",
         243 => x"232ef107",
         244 => x"f3272034",
         245 => x"1307b000",
         246 => x"6388e708",
         247 => x"13073000",
         248 => x"638ce70e",
         249 => x"03258102",
         250 => x"832fc107",
         251 => x"032f8107",
         252 => x"832e4107",
         253 => x"032e0107",
         254 => x"832dc106",
         255 => x"032d8106",
         256 => x"832c4106",
         257 => x"032c0106",
         258 => x"832bc105",
         259 => x"032b8105",
         260 => x"832a4105",
         261 => x"032a0105",
         262 => x"8329c104",
         263 => x"03298104",
         264 => x"83284104",
         265 => x"03280104",
         266 => x"8327c103",
         267 => x"03278103",
         268 => x"83264103",
         269 => x"03260103",
         270 => x"8325c102",
         271 => x"83244102",
         272 => x"03240102",
         273 => x"8323c101",
         274 => x"03238101",
         275 => x"83224101",
         276 => x"03220101",
         277 => x"8321c100",
         278 => x"03218100",
         279 => x"83204100",
         280 => x"13010108",
         281 => x"73002030",
         282 => x"9307600d",
         283 => x"638ef806",
         284 => x"9307900a",
         285 => x"6382f818",
         286 => x"63c41703",
         287 => x"938878fc",
         288 => x"93074002",
         289 => x"63e0170b",
         290 => x"b7370000",
         291 => x"93874700",
         292 => x"93982800",
         293 => x"b388f800",
         294 => x"83a70800",
         295 => x"67800700",
         296 => x"938808c0",
         297 => x"9307f000",
         298 => x"63ee1707",
         299 => x"b7370000",
         300 => x"93878709",
         301 => x"93982800",
         302 => x"b388f800",
         303 => x"83a70800",
         304 => x"67800700",
         305 => x"b7270000",
         306 => x"23a2f500",
         307 => x"93070000",
         308 => x"13850700",
         309 => x"6ff05ff1",
         310 => x"13050100",
         311 => x"ef004018",
         312 => x"03258102",
         313 => x"6ff05ff0",
         314 => x"63180500",
         315 => x"13858189",
         316 => x"13050500",
         317 => x"6ff05fef",
         318 => x"b7870020",
         319 => x"93870700",
         320 => x"13070040",
         321 => x"b387e740",
         322 => x"e364f5fe",
         323 => x"ef10005b",
         324 => x"9307c000",
         325 => x"2320f500",
         326 => x"1305f0ff",
         327 => x"13050500",
         328 => x"6ff09fec",
         329 => x"ef108059",
         330 => x"93078005",
         331 => x"2320f500",
         332 => x"9307f0ff",
         333 => x"13850700",
         334 => x"6ff01feb",
         335 => x"ef100058",
         336 => x"93079000",
         337 => x"2320f500",
         338 => x"9307f0ff",
         339 => x"13850700",
         340 => x"6ff09fe9",
         341 => x"93070000",
         342 => x"13850700",
         343 => x"6ff0dfe8",
         344 => x"ef10c055",
         345 => x"9307d000",
         346 => x"2320f500",
         347 => x"9307f0ff",
         348 => x"13850700",
         349 => x"6ff05fe7",
         350 => x"ef104054",
         351 => x"9307f001",
         352 => x"2320f500",
         353 => x"9307f0ff",
         354 => x"13850700",
         355 => x"6ff0dfe5",
         356 => x"ef10c052",
         357 => x"93072000",
         358 => x"2320f500",
         359 => x"9307f0ff",
         360 => x"13850700",
         361 => x"6ff05fe4",
         362 => x"13090600",
         363 => x"13840500",
         364 => x"635cc000",
         365 => x"b384c500",
         366 => x"eff0dfce",
         367 => x"2300a400",
         368 => x"13041400",
         369 => x"e31a94fe",
         370 => x"13050900",
         371 => x"6ff0dfe1",
         372 => x"13090600",
         373 => x"13840500",
         374 => x"e358c0fe",
         375 => x"b384c500",
         376 => x"03450400",
         377 => x"13041400",
         378 => x"eff09fc9",
         379 => x"e39a84fe",
         380 => x"13050900",
         381 => x"6ff05fdf",
         382 => x"13090000",
         383 => x"93040500",
         384 => x"13040900",
         385 => x"93090900",
         386 => x"93070900",
         387 => x"732410c8",
         388 => x"f32910c0",
         389 => x"f32710c8",
         390 => x"e31af4fe",
         391 => x"37460f00",
         392 => x"13060624",
         393 => x"93060000",
         394 => x"13850900",
         395 => x"93050400",
         396 => x"ef005068",
         397 => x"37460f00",
         398 => x"23a4a400",
         399 => x"13060624",
         400 => x"93060000",
         401 => x"13850900",
         402 => x"93050400",
         403 => x"ef009023",
         404 => x"23a0a400",
         405 => x"23a2b400",
         406 => x"13050900",
         407 => x"6ff0dfd8",
         408 => x"37350000",
         409 => x"130101ff",
         410 => x"1305052d",
         411 => x"23261100",
         412 => x"23248100",
         413 => x"23229100",
         414 => x"23202101",
         415 => x"eff09fa3",
         416 => x"73294034",
         417 => x"93040002",
         418 => x"37040080",
         419 => x"33758900",
         420 => x"3335a000",
         421 => x"13050503",
         422 => x"9384f4ff",
         423 => x"eff09f9f",
         424 => x"13541400",
         425 => x"e39404fe",
         426 => x"03248100",
         427 => x"8320c100",
         428 => x"83244100",
         429 => x"03290100",
         430 => x"37350000",
         431 => x"13054520",
         432 => x"13010101",
         433 => x"6ff01f9f",
         434 => x"130101ff",
         435 => x"2322f100",
         436 => x"b70700f0",
         437 => x"2324e100",
         438 => x"03a74708",
         439 => x"2326d100",
         440 => x"8326c100",
         441 => x"1377f7fe",
         442 => x"23a2e708",
         443 => x"03a74700",
         444 => x"13471700",
         445 => x"23a2e700",
         446 => x"03278100",
         447 => x"83274100",
         448 => x"13010101",
         449 => x"73002030",
         450 => x"6f000000",
         451 => x"130101fe",
         452 => x"2326f100",
         453 => x"b70700f0",
         454 => x"232eb100",
         455 => x"2328e100",
         456 => x"83a5470f",
         457 => x"03a7070f",
         458 => x"232ad100",
         459 => x"b7860100",
         460 => x"232cc100",
         461 => x"9386066a",
         462 => x"1306f0ff",
         463 => x"23aec70e",
         464 => x"b306d700",
         465 => x"23acc70e",
         466 => x"33b7e600",
         467 => x"23acd70e",
         468 => x"3307b700",
         469 => x"23aee70e",
         470 => x"03a74700",
         471 => x"8325c101",
         472 => x"03268101",
         473 => x"13472700",
         474 => x"23a2e700",
         475 => x"83264101",
         476 => x"03270101",
         477 => x"8327c100",
         478 => x"13010102",
         479 => x"73002030",
         480 => x"130101ff",
         481 => x"2326e100",
         482 => x"370700f0",
         483 => x"2324f100",
         484 => x"8327c702",
         485 => x"93f74700",
         486 => x"638a0700",
         487 => x"83274700",
         488 => x"93c74700",
         489 => x"2322f700",
         490 => x"83270702",
         491 => x"0327c100",
         492 => x"83278100",
         493 => x"13010101",
         494 => x"73002030",
         495 => x"13030500",
         496 => x"138e0500",
         497 => x"93080000",
         498 => x"63dc0500",
         499 => x"b337a000",
         500 => x"330eb040",
         501 => x"330efe40",
         502 => x"3303a040",
         503 => x"9308f0ff",
         504 => x"63dc0600",
         505 => x"b337c000",
         506 => x"b306d040",
         507 => x"93c8f8ff",
         508 => x"b386f640",
         509 => x"3306c040",
         510 => x"13070600",
         511 => x"13080300",
         512 => x"93070e00",
         513 => x"639c0628",
         514 => x"b7350000",
         515 => x"9385850d",
         516 => x"6376ce0e",
         517 => x"b7060100",
         518 => x"6378d60c",
         519 => x"93360610",
         520 => x"93c61600",
         521 => x"93963600",
         522 => x"3355d600",
         523 => x"b385a500",
         524 => x"83c50500",
         525 => x"13050002",
         526 => x"b386d500",
         527 => x"b305d540",
         528 => x"630cd500",
         529 => x"b317be00",
         530 => x"b356d300",
         531 => x"3317b600",
         532 => x"b3e7f600",
         533 => x"3318b300",
         534 => x"93550701",
         535 => x"33deb702",
         536 => x"13160701",
         537 => x"13560601",
         538 => x"b3f7b702",
         539 => x"13050e00",
         540 => x"3303c603",
         541 => x"93960701",
         542 => x"93570801",
         543 => x"b3e7d700",
         544 => x"63fe6700",
         545 => x"b387e700",
         546 => x"1305feff",
         547 => x"63e8e700",
         548 => x"63f66700",
         549 => x"1305eeff",
         550 => x"b387e700",
         551 => x"b3876740",
         552 => x"33d3b702",
         553 => x"13180801",
         554 => x"13580801",
         555 => x"b3f7b702",
         556 => x"b3066602",
         557 => x"93970701",
         558 => x"3368f800",
         559 => x"93070300",
         560 => x"637cd800",
         561 => x"33080701",
         562 => x"9307f3ff",
         563 => x"6366e800",
         564 => x"6374d800",
         565 => x"9307e3ff",
         566 => x"13150501",
         567 => x"3365f500",
         568 => x"93050000",
         569 => x"6f00000e",
         570 => x"37050001",
         571 => x"93060001",
         572 => x"e36ca6f2",
         573 => x"93068001",
         574 => x"6ff01ff3",
         575 => x"63140600",
         576 => x"73001000",
         577 => x"b7070100",
         578 => x"637af60c",
         579 => x"93360610",
         580 => x"93c61600",
         581 => x"93963600",
         582 => x"b357d600",
         583 => x"b385f500",
         584 => x"83c70500",
         585 => x"b387d700",
         586 => x"93060002",
         587 => x"b385f640",
         588 => x"6390f60c",
         589 => x"b307ce40",
         590 => x"93051000",
         591 => x"13530701",
         592 => x"b3de6702",
         593 => x"13160701",
         594 => x"13560601",
         595 => x"93560801",
         596 => x"b3f76702",
         597 => x"13850e00",
         598 => x"330ed603",
         599 => x"93970701",
         600 => x"b3e7f600",
         601 => x"63fec701",
         602 => x"b387e700",
         603 => x"1385feff",
         604 => x"63e8e700",
         605 => x"63f6c701",
         606 => x"1385eeff",
         607 => x"b387e700",
         608 => x"b387c741",
         609 => x"33de6702",
         610 => x"13180801",
         611 => x"13580801",
         612 => x"b3f76702",
         613 => x"b306c603",
         614 => x"93970701",
         615 => x"3368f800",
         616 => x"93070e00",
         617 => x"637cd800",
         618 => x"33080701",
         619 => x"9307feff",
         620 => x"6366e800",
         621 => x"6374d800",
         622 => x"9307eeff",
         623 => x"13150501",
         624 => x"3365f500",
         625 => x"638a0800",
         626 => x"b337a000",
         627 => x"b305b040",
         628 => x"b385f540",
         629 => x"3305a040",
         630 => x"67800000",
         631 => x"b7070001",
         632 => x"93060001",
         633 => x"e36af6f2",
         634 => x"93068001",
         635 => x"6ff0dff2",
         636 => x"3317b600",
         637 => x"b356fe00",
         638 => x"13550701",
         639 => x"331ebe00",
         640 => x"b357f300",
         641 => x"b3e7c701",
         642 => x"33dea602",
         643 => x"13160701",
         644 => x"13560601",
         645 => x"3318b300",
         646 => x"b3f6a602",
         647 => x"3303c603",
         648 => x"93950601",
         649 => x"93d60701",
         650 => x"b3e6b600",
         651 => x"93050e00",
         652 => x"63fe6600",
         653 => x"b386e600",
         654 => x"9305feff",
         655 => x"63e8e600",
         656 => x"63f66600",
         657 => x"9305eeff",
         658 => x"b386e600",
         659 => x"b3866640",
         660 => x"33d3a602",
         661 => x"93970701",
         662 => x"93d70701",
         663 => x"b3f6a602",
         664 => x"33066602",
         665 => x"93960601",
         666 => x"b3e7d700",
         667 => x"93060300",
         668 => x"63fec700",
         669 => x"b387e700",
         670 => x"9306f3ff",
         671 => x"63e8e700",
         672 => x"63f6c700",
         673 => x"9306e3ff",
         674 => x"b387e700",
         675 => x"93950501",
         676 => x"b387c740",
         677 => x"b3e5d500",
         678 => x"6ff05fea",
         679 => x"6366de18",
         680 => x"b7070100",
         681 => x"63f4f604",
         682 => x"13b70610",
         683 => x"13471700",
         684 => x"13173700",
         685 => x"b7370000",
         686 => x"b3d5e600",
         687 => x"9387870d",
         688 => x"b387b700",
         689 => x"83c70700",
         690 => x"b387e700",
         691 => x"13070002",
         692 => x"b305f740",
         693 => x"6316f702",
         694 => x"13051000",
         695 => x"e3e4c6ef",
         696 => x"3335c300",
         697 => x"13451500",
         698 => x"6ff0dfed",
         699 => x"b7070001",
         700 => x"13070001",
         701 => x"e3e0f6fc",
         702 => x"13078001",
         703 => x"6ff09ffb",
         704 => x"3357f600",
         705 => x"b396b600",
         706 => x"b366d700",
         707 => x"3357fe00",
         708 => x"331ebe00",
         709 => x"b357f300",
         710 => x"b3e7c701",
         711 => x"13de0601",
         712 => x"335fc703",
         713 => x"13980601",
         714 => x"13580801",
         715 => x"3316b600",
         716 => x"3377c703",
         717 => x"b30ee803",
         718 => x"13150701",
         719 => x"13d70701",
         720 => x"3367a700",
         721 => x"13050f00",
         722 => x"637ed701",
         723 => x"3307d700",
         724 => x"1305ffff",
         725 => x"6368d700",
         726 => x"6376d701",
         727 => x"1305efff",
         728 => x"3307d700",
         729 => x"3307d741",
         730 => x"b35ec703",
         731 => x"93970701",
         732 => x"93d70701",
         733 => x"3377c703",
         734 => x"3308d803",
         735 => x"13170701",
         736 => x"b3e7e700",
         737 => x"13870e00",
         738 => x"63fe0701",
         739 => x"b387d700",
         740 => x"1387feff",
         741 => x"63e8d700",
         742 => x"63f60701",
         743 => x"1387eeff",
         744 => x"b387d700",
         745 => x"13150501",
         746 => x"b70e0100",
         747 => x"3365e500",
         748 => x"9386feff",
         749 => x"3377d500",
         750 => x"b3870741",
         751 => x"b376d600",
         752 => x"13580501",
         753 => x"13560601",
         754 => x"330ed702",
         755 => x"b306d802",
         756 => x"3307c702",
         757 => x"3308c802",
         758 => x"3306d700",
         759 => x"13570e01",
         760 => x"3307c700",
         761 => x"6374d700",
         762 => x"3308d801",
         763 => x"93560701",
         764 => x"b3860601",
         765 => x"63e6d702",
         766 => x"e394d7ce",
         767 => x"b7070100",
         768 => x"9387f7ff",
         769 => x"3377f700",
         770 => x"13170701",
         771 => x"337efe00",
         772 => x"3313b300",
         773 => x"3307c701",
         774 => x"93050000",
         775 => x"e374e3da",
         776 => x"1305f5ff",
         777 => x"6ff0dfcb",
         778 => x"93050000",
         779 => x"13050000",
         780 => x"6ff05fd9",
         781 => x"138e0500",
         782 => x"13080000",
         783 => x"63dc0500",
         784 => x"b337a000",
         785 => x"b305b040",
         786 => x"338ef540",
         787 => x"3305a040",
         788 => x"1308f0ff",
         789 => x"63da0600",
         790 => x"b337c000",
         791 => x"b306d040",
         792 => x"b386f640",
         793 => x"3306c040",
         794 => x"93080600",
         795 => x"93070500",
         796 => x"93050e00",
         797 => x"63940624",
         798 => x"37370000",
         799 => x"1307870d",
         800 => x"6376ce0e",
         801 => x"b7060100",
         802 => x"6378d60c",
         803 => x"93360610",
         804 => x"93c61600",
         805 => x"93963600",
         806 => x"3353d600",
         807 => x"33076700",
         808 => x"03470700",
         809 => x"3307d700",
         810 => x"93060002",
         811 => x"3383e640",
         812 => x"638ce600",
         813 => x"b3156e00",
         814 => x"3357e500",
         815 => x"b3186600",
         816 => x"b365b700",
         817 => x"b3176500",
         818 => x"93d60801",
         819 => x"33d7d502",
         820 => x"13950801",
         821 => x"13550501",
         822 => x"b3f5d502",
         823 => x"3307a702",
         824 => x"13960501",
         825 => x"93d50701",
         826 => x"b3e5c500",
         827 => x"63fae500",
         828 => x"b3851501",
         829 => x"63e61501",
         830 => x"63f4e500",
         831 => x"b3851501",
         832 => x"b385e540",
         833 => x"33d7d502",
         834 => x"93970701",
         835 => x"93d70701",
         836 => x"b3f5d502",
         837 => x"3307a702",
         838 => x"93950501",
         839 => x"b3e7b700",
         840 => x"63fae700",
         841 => x"b3871701",
         842 => x"63e61701",
         843 => x"63f4e700",
         844 => x"b3871701",
         845 => x"b387e740",
         846 => x"33d56700",
         847 => x"93050000",
         848 => x"630a0800",
         849 => x"b337a000",
         850 => x"b305b040",
         851 => x"b385f540",
         852 => x"3305a040",
         853 => x"67800000",
         854 => x"37030001",
         855 => x"93060001",
         856 => x"e36c66f2",
         857 => x"93068001",
         858 => x"6ff01ff3",
         859 => x"63140600",
         860 => x"73001000",
         861 => x"b7060100",
         862 => x"6372d60a",
         863 => x"93360610",
         864 => x"93c61600",
         865 => x"93963600",
         866 => x"b355d600",
         867 => x"3307b700",
         868 => x"03470700",
         869 => x"3307d700",
         870 => x"93060002",
         871 => x"3383e640",
         872 => x"6398e608",
         873 => x"3307ce40",
         874 => x"93d50801",
         875 => x"3356b702",
         876 => x"13950801",
         877 => x"13550501",
         878 => x"93d60701",
         879 => x"3377b702",
         880 => x"3306a602",
         881 => x"13170701",
         882 => x"33e7e600",
         883 => x"637ac700",
         884 => x"33071701",
         885 => x"63661701",
         886 => x"6374c700",
         887 => x"33071701",
         888 => x"3307c740",
         889 => x"b356b702",
         890 => x"93970701",
         891 => x"93d70701",
         892 => x"3377b702",
         893 => x"b386a602",
         894 => x"13170701",
         895 => x"b3e7e700",
         896 => x"63fad700",
         897 => x"b3871701",
         898 => x"63e61701",
         899 => x"63f4d700",
         900 => x"b3871701",
         901 => x"b387d740",
         902 => x"6ff01ff2",
         903 => x"b7050001",
         904 => x"93060001",
         905 => x"e362b6f6",
         906 => x"93068001",
         907 => x"6ff0dff5",
         908 => x"b3186600",
         909 => x"b356ee00",
         910 => x"b3156e00",
         911 => x"3357e500",
         912 => x"b3176500",
         913 => x"13d50801",
         914 => x"3367b700",
         915 => x"b3d5a602",
         916 => x"139e0801",
         917 => x"135e0e01",
         918 => x"b3f6a602",
         919 => x"b385c503",
         920 => x"13960601",
         921 => x"93560701",
         922 => x"b3e6c600",
         923 => x"63fab600",
         924 => x"b3861601",
         925 => x"63e61601",
         926 => x"63f4b600",
         927 => x"b3861601",
         928 => x"b386b640",
         929 => x"33d6a602",
         930 => x"13170701",
         931 => x"13570701",
         932 => x"b3f6a602",
         933 => x"3306c603",
         934 => x"93960601",
         935 => x"3367d700",
         936 => x"637ac700",
         937 => x"33071701",
         938 => x"63661701",
         939 => x"6374c700",
         940 => x"33071701",
         941 => x"3307c740",
         942 => x"6ff01fef",
         943 => x"e362dee8",
         944 => x"37070100",
         945 => x"63fce604",
         946 => x"13b70610",
         947 => x"13471700",
         948 => x"13173700",
         949 => x"b7380000",
         950 => x"33d3e600",
         951 => x"9388880d",
         952 => x"b3886800",
         953 => x"03c30800",
         954 => x"3303e300",
         955 => x"13070002",
         956 => x"b3086740",
         957 => x"631e6702",
         958 => x"63e4c601",
         959 => x"636cc500",
         960 => x"3306c540",
         961 => x"b306de40",
         962 => x"b335c500",
         963 => x"b385b640",
         964 => x"93070600",
         965 => x"13850700",
         966 => x"6ff09fe2",
         967 => x"b7080001",
         968 => x"13070001",
         969 => x"e3e816fb",
         970 => x"13078001",
         971 => x"6ff09ffa",
         972 => x"b3576600",
         973 => x"b3961601",
         974 => x"b3e6d700",
         975 => x"33576e00",
         976 => x"93de0601",
         977 => x"b35fd703",
         978 => x"b3151e01",
         979 => x"139e0601",
         980 => x"135e0e01",
         981 => x"b3576500",
         982 => x"b3e5b700",
         983 => x"93d70501",
         984 => x"33161601",
         985 => x"33151501",
         986 => x"3377d703",
         987 => x"330ffe03",
         988 => x"13170701",
         989 => x"b3e7e700",
         990 => x"13870f00",
         991 => x"63fee701",
         992 => x"b387d700",
         993 => x"1387ffff",
         994 => x"63e8d700",
         995 => x"63f6e701",
         996 => x"1387efff",
         997 => x"b387d700",
         998 => x"b387e741",
         999 => x"33dfd703",
        1000 => x"93950501",
        1001 => x"93d50501",
        1002 => x"b3f7d703",
        1003 => x"330eee03",
        1004 => x"93970701",
        1005 => x"b3e5f500",
        1006 => x"93070f00",
        1007 => x"63fec501",
        1008 => x"b385d500",
        1009 => x"9307ffff",
        1010 => x"63e8d500",
        1011 => x"63f6c501",
        1012 => x"9307efff",
        1013 => x"b385d500",
        1014 => x"13170701",
        1015 => x"b70f0100",
        1016 => x"3367f700",
        1017 => x"b385c541",
        1018 => x"138effff",
        1019 => x"b377c701",
        1020 => x"935e0601",
        1021 => x"13570701",
        1022 => x"337ec601",
        1023 => x"338fc703",
        1024 => x"330ec703",
        1025 => x"b387d703",
        1026 => x"3307d703",
        1027 => x"b38ec701",
        1028 => x"93570f01",
        1029 => x"b387d701",
        1030 => x"63f4c701",
        1031 => x"3307f701",
        1032 => x"13de0701",
        1033 => x"3307ee00",
        1034 => x"370e0100",
        1035 => x"130efeff",
        1036 => x"b3f7c701",
        1037 => x"93970701",
        1038 => x"337fcf01",
        1039 => x"b387e701",
        1040 => x"63e6e500",
        1041 => x"639ee500",
        1042 => x"637cf500",
        1043 => x"3386c740",
        1044 => x"b3b7c700",
        1045 => x"b387d700",
        1046 => x"3307f740",
        1047 => x"93070600",
        1048 => x"b307f540",
        1049 => x"3335f500",
        1050 => x"b385e540",
        1051 => x"b385a540",
        1052 => x"33936500",
        1053 => x"b3d71701",
        1054 => x"3365f300",
        1055 => x"b3d51501",
        1056 => x"6ff01fcc",
        1057 => x"13030500",
        1058 => x"93880500",
        1059 => x"13070600",
        1060 => x"13080500",
        1061 => x"93870500",
        1062 => x"63920628",
        1063 => x"b7350000",
        1064 => x"9385850d",
        1065 => x"63f6c80e",
        1066 => x"b7060100",
        1067 => x"6378d60c",
        1068 => x"93360610",
        1069 => x"93c61600",
        1070 => x"93963600",
        1071 => x"3355d600",
        1072 => x"b385a500",
        1073 => x"83c50500",
        1074 => x"13050002",
        1075 => x"b386d500",
        1076 => x"b305d540",
        1077 => x"630cd500",
        1078 => x"b397b800",
        1079 => x"b356d300",
        1080 => x"3317b600",
        1081 => x"b3e7f600",
        1082 => x"3318b300",
        1083 => x"93550701",
        1084 => x"33d3b702",
        1085 => x"13160701",
        1086 => x"13560601",
        1087 => x"b3f7b702",
        1088 => x"13050300",
        1089 => x"b3086602",
        1090 => x"93960701",
        1091 => x"93570801",
        1092 => x"b3e7d700",
        1093 => x"63fe1701",
        1094 => x"b387e700",
        1095 => x"1305f3ff",
        1096 => x"63e8e700",
        1097 => x"63f61701",
        1098 => x"1305e3ff",
        1099 => x"b387e700",
        1100 => x"b3871741",
        1101 => x"b3d8b702",
        1102 => x"13180801",
        1103 => x"13580801",
        1104 => x"b3f7b702",
        1105 => x"b3061603",
        1106 => x"93970701",
        1107 => x"3368f800",
        1108 => x"93870800",
        1109 => x"637cd800",
        1110 => x"33080701",
        1111 => x"9387f8ff",
        1112 => x"6366e800",
        1113 => x"6374d800",
        1114 => x"9387e8ff",
        1115 => x"13150501",
        1116 => x"3365f500",
        1117 => x"93050000",
        1118 => x"67800000",
        1119 => x"37050001",
        1120 => x"93060001",
        1121 => x"e36ca6f2",
        1122 => x"93068001",
        1123 => x"6ff01ff3",
        1124 => x"63140600",
        1125 => x"73001000",
        1126 => x"b7070100",
        1127 => x"6370f60c",
        1128 => x"93360610",
        1129 => x"93c61600",
        1130 => x"93963600",
        1131 => x"b357d600",
        1132 => x"b385f500",
        1133 => x"83c70500",
        1134 => x"b387d700",
        1135 => x"93060002",
        1136 => x"b385f640",
        1137 => x"6396f60a",
        1138 => x"b387c840",
        1139 => x"93051000",
        1140 => x"93580701",
        1141 => x"33de1703",
        1142 => x"13160701",
        1143 => x"13560601",
        1144 => x"93560801",
        1145 => x"b3f71703",
        1146 => x"13050e00",
        1147 => x"3303c603",
        1148 => x"93970701",
        1149 => x"b3e7f600",
        1150 => x"63fe6700",
        1151 => x"b387e700",
        1152 => x"1305feff",
        1153 => x"63e8e700",
        1154 => x"63f66700",
        1155 => x"1305eeff",
        1156 => x"b387e700",
        1157 => x"b3876740",
        1158 => x"33d31703",
        1159 => x"13180801",
        1160 => x"13580801",
        1161 => x"b3f71703",
        1162 => x"b3066602",
        1163 => x"93970701",
        1164 => x"3368f800",
        1165 => x"93070300",
        1166 => x"637cd800",
        1167 => x"33080701",
        1168 => x"9307f3ff",
        1169 => x"6366e800",
        1170 => x"6374d800",
        1171 => x"9307e3ff",
        1172 => x"13150501",
        1173 => x"3365f500",
        1174 => x"67800000",
        1175 => x"b7070001",
        1176 => x"93060001",
        1177 => x"e364f6f4",
        1178 => x"93068001",
        1179 => x"6ff01ff4",
        1180 => x"3317b600",
        1181 => x"b3d6f800",
        1182 => x"13550701",
        1183 => x"b357f300",
        1184 => x"3318b300",
        1185 => x"33d3a602",
        1186 => x"13160701",
        1187 => x"b398b800",
        1188 => x"13560601",
        1189 => x"b3e71701",
        1190 => x"b3f6a602",
        1191 => x"b3086602",
        1192 => x"93950601",
        1193 => x"93d60701",
        1194 => x"b3e6b600",
        1195 => x"93050300",
        1196 => x"63fe1601",
        1197 => x"b386e600",
        1198 => x"9305f3ff",
        1199 => x"63e8e600",
        1200 => x"63f61601",
        1201 => x"9305e3ff",
        1202 => x"b386e600",
        1203 => x"b3861641",
        1204 => x"b3d8a602",
        1205 => x"93970701",
        1206 => x"93d70701",
        1207 => x"b3f6a602",
        1208 => x"33061603",
        1209 => x"93960601",
        1210 => x"b3e7d700",
        1211 => x"93860800",
        1212 => x"63fec700",
        1213 => x"b387e700",
        1214 => x"9386f8ff",
        1215 => x"63e8e700",
        1216 => x"63f6c700",
        1217 => x"9386e8ff",
        1218 => x"b387e700",
        1219 => x"93950501",
        1220 => x"b387c740",
        1221 => x"b3e5d500",
        1222 => x"6ff09feb",
        1223 => x"63e6d518",
        1224 => x"b7070100",
        1225 => x"63f4f604",
        1226 => x"13b70610",
        1227 => x"13471700",
        1228 => x"13173700",
        1229 => x"b7370000",
        1230 => x"b3d5e600",
        1231 => x"9387870d",
        1232 => x"b387b700",
        1233 => x"83c70700",
        1234 => x"b387e700",
        1235 => x"13070002",
        1236 => x"b305f740",
        1237 => x"6316f702",
        1238 => x"13051000",
        1239 => x"e3ee16e1",
        1240 => x"3335c300",
        1241 => x"13451500",
        1242 => x"67800000",
        1243 => x"b7070001",
        1244 => x"13070001",
        1245 => x"e3e0f6fc",
        1246 => x"13078001",
        1247 => x"6ff09ffb",
        1248 => x"3357f600",
        1249 => x"b396b600",
        1250 => x"b366d700",
        1251 => x"33d7f800",
        1252 => x"b398b800",
        1253 => x"b357f300",
        1254 => x"b3e71701",
        1255 => x"93d80601",
        1256 => x"b35e1703",
        1257 => x"13980601",
        1258 => x"13580801",
        1259 => x"3316b600",
        1260 => x"33771703",
        1261 => x"330ed803",
        1262 => x"13150701",
        1263 => x"13d70701",
        1264 => x"3367a700",
        1265 => x"13850e00",
        1266 => x"637ec701",
        1267 => x"3307d700",
        1268 => x"1385feff",
        1269 => x"6368d700",
        1270 => x"6376c701",
        1271 => x"1385eeff",
        1272 => x"3307d700",
        1273 => x"3307c741",
        1274 => x"335e1703",
        1275 => x"93970701",
        1276 => x"93d70701",
        1277 => x"33771703",
        1278 => x"3308c803",
        1279 => x"13170701",
        1280 => x"b3e7e700",
        1281 => x"13070e00",
        1282 => x"63fe0701",
        1283 => x"b387d700",
        1284 => x"1307feff",
        1285 => x"63e8d700",
        1286 => x"63f60701",
        1287 => x"1307eeff",
        1288 => x"b387d700",
        1289 => x"13150501",
        1290 => x"370e0100",
        1291 => x"3365e500",
        1292 => x"9306feff",
        1293 => x"3377d500",
        1294 => x"b3870741",
        1295 => x"b376d600",
        1296 => x"13580501",
        1297 => x"13560601",
        1298 => x"b308d702",
        1299 => x"b306d802",
        1300 => x"3307c702",
        1301 => x"3308c802",
        1302 => x"3306d700",
        1303 => x"13d70801",
        1304 => x"3307c700",
        1305 => x"6374d700",
        1306 => x"3308c801",
        1307 => x"93560701",
        1308 => x"b3860601",
        1309 => x"63e6d702",
        1310 => x"e39ed7ce",
        1311 => x"b7070100",
        1312 => x"9387f7ff",
        1313 => x"3377f700",
        1314 => x"13170701",
        1315 => x"b3f8f800",
        1316 => x"3313b300",
        1317 => x"33071701",
        1318 => x"93050000",
        1319 => x"e37ee3cc",
        1320 => x"1305f5ff",
        1321 => x"6ff01fcd",
        1322 => x"93050000",
        1323 => x"13050000",
        1324 => x"67800000",
        1325 => x"13080600",
        1326 => x"93070500",
        1327 => x"13870500",
        1328 => x"63960620",
        1329 => x"b7380000",
        1330 => x"9388880d",
        1331 => x"63fcc50c",
        1332 => x"b7060100",
        1333 => x"637ed60a",
        1334 => x"93360610",
        1335 => x"93c61600",
        1336 => x"93963600",
        1337 => x"3353d600",
        1338 => x"b3886800",
        1339 => x"83c80800",
        1340 => x"13030002",
        1341 => x"b386d800",
        1342 => x"b308d340",
        1343 => x"630cd300",
        1344 => x"33971501",
        1345 => x"b356d500",
        1346 => x"33181601",
        1347 => x"33e7e600",
        1348 => x"b3171501",
        1349 => x"13560801",
        1350 => x"b356c702",
        1351 => x"13150801",
        1352 => x"13550501",
        1353 => x"3377c702",
        1354 => x"b386a602",
        1355 => x"93150701",
        1356 => x"13d70701",
        1357 => x"3367b700",
        1358 => x"637ad700",
        1359 => x"33070701",
        1360 => x"63660701",
        1361 => x"6374d700",
        1362 => x"33070701",
        1363 => x"3307d740",
        1364 => x"b356c702",
        1365 => x"3377c702",
        1366 => x"b386a602",
        1367 => x"93970701",
        1368 => x"13170701",
        1369 => x"93d70701",
        1370 => x"b3e7e700",
        1371 => x"63fad700",
        1372 => x"b3870701",
        1373 => x"63e60701",
        1374 => x"63f4d700",
        1375 => x"b3870701",
        1376 => x"b387d740",
        1377 => x"33d51701",
        1378 => x"93050000",
        1379 => x"67800000",
        1380 => x"37030001",
        1381 => x"93060001",
        1382 => x"e36666f4",
        1383 => x"93068001",
        1384 => x"6ff05ff4",
        1385 => x"63140600",
        1386 => x"73001000",
        1387 => x"37070100",
        1388 => x"637ee606",
        1389 => x"93360610",
        1390 => x"93c61600",
        1391 => x"93963600",
        1392 => x"3357d600",
        1393 => x"b388e800",
        1394 => x"03c70800",
        1395 => x"3307d700",
        1396 => x"93060002",
        1397 => x"b388e640",
        1398 => x"6394e606",
        1399 => x"3387c540",
        1400 => x"93550801",
        1401 => x"3356b702",
        1402 => x"13150801",
        1403 => x"13550501",
        1404 => x"93d60701",
        1405 => x"3377b702",
        1406 => x"3306a602",
        1407 => x"13170701",
        1408 => x"33e7e600",
        1409 => x"637ac700",
        1410 => x"33070701",
        1411 => x"63660701",
        1412 => x"6374c700",
        1413 => x"33070701",
        1414 => x"3307c740",
        1415 => x"b356b702",
        1416 => x"3377b702",
        1417 => x"b386a602",
        1418 => x"6ff05ff3",
        1419 => x"37070001",
        1420 => x"93060001",
        1421 => x"e366e6f8",
        1422 => x"93068001",
        1423 => x"6ff05ff8",
        1424 => x"33181601",
        1425 => x"b3d6e500",
        1426 => x"b3171501",
        1427 => x"b3951501",
        1428 => x"3357e500",
        1429 => x"13550801",
        1430 => x"3367b700",
        1431 => x"b3d5a602",
        1432 => x"13130801",
        1433 => x"13530301",
        1434 => x"b3f6a602",
        1435 => x"b3856502",
        1436 => x"13960601",
        1437 => x"93560701",
        1438 => x"b3e6c600",
        1439 => x"63fab600",
        1440 => x"b3860601",
        1441 => x"63e60601",
        1442 => x"63f4b600",
        1443 => x"b3860601",
        1444 => x"b386b640",
        1445 => x"33d6a602",
        1446 => x"13170701",
        1447 => x"13570701",
        1448 => x"b3f6a602",
        1449 => x"33066602",
        1450 => x"93960601",
        1451 => x"3367d700",
        1452 => x"637ac700",
        1453 => x"33070701",
        1454 => x"63660701",
        1455 => x"6374c700",
        1456 => x"33070701",
        1457 => x"3307c740",
        1458 => x"6ff09ff1",
        1459 => x"63e4d51c",
        1460 => x"37080100",
        1461 => x"63fe0605",
        1462 => x"13b80610",
        1463 => x"13481800",
        1464 => x"13183800",
        1465 => x"b7380000",
        1466 => x"33d30601",
        1467 => x"9388880d",
        1468 => x"b3886800",
        1469 => x"83c80800",
        1470 => x"13030002",
        1471 => x"b3880801",
        1472 => x"33081341",
        1473 => x"63101305",
        1474 => x"63e4b600",
        1475 => x"636cc500",
        1476 => x"3306c540",
        1477 => x"b386d540",
        1478 => x"3337c500",
        1479 => x"3387e640",
        1480 => x"93070600",
        1481 => x"13850700",
        1482 => x"93050700",
        1483 => x"67800000",
        1484 => x"b7080001",
        1485 => x"13080001",
        1486 => x"e3e616fb",
        1487 => x"13088001",
        1488 => x"6ff05ffa",
        1489 => x"b3960601",
        1490 => x"33531601",
        1491 => x"3363d300",
        1492 => x"135e0301",
        1493 => x"b3d61501",
        1494 => x"33dfc603",
        1495 => x"13170301",
        1496 => x"13570701",
        1497 => x"b3970501",
        1498 => x"b3551501",
        1499 => x"b3e5f500",
        1500 => x"93d70501",
        1501 => x"33160601",
        1502 => x"33150501",
        1503 => x"b3f6c603",
        1504 => x"b30ee703",
        1505 => x"93960601",
        1506 => x"b3e7d700",
        1507 => x"93060f00",
        1508 => x"63fed701",
        1509 => x"b3876700",
        1510 => x"9306ffff",
        1511 => x"63e86700",
        1512 => x"63f6d701",
        1513 => x"9306efff",
        1514 => x"b3876700",
        1515 => x"b387d741",
        1516 => x"b3dec703",
        1517 => x"93950501",
        1518 => x"93d50501",
        1519 => x"b3f7c703",
        1520 => x"3307d703",
        1521 => x"93970701",
        1522 => x"b3e5f500",
        1523 => x"93870e00",
        1524 => x"63fee500",
        1525 => x"b3856500",
        1526 => x"9387feff",
        1527 => x"63e86500",
        1528 => x"63f6e500",
        1529 => x"9387eeff",
        1530 => x"b3856500",
        1531 => x"93960601",
        1532 => x"370f0100",
        1533 => x"b3e6f600",
        1534 => x"9307ffff",
        1535 => x"135e0601",
        1536 => x"b385e540",
        1537 => x"33f7f600",
        1538 => x"93d60601",
        1539 => x"b377f600",
        1540 => x"b30ef702",
        1541 => x"b387f602",
        1542 => x"3307c703",
        1543 => x"b386c603",
        1544 => x"330ef700",
        1545 => x"13d70e01",
        1546 => x"3307c701",
        1547 => x"6374f700",
        1548 => x"b386e601",
        1549 => x"93570701",
        1550 => x"b387d700",
        1551 => x"b7060100",
        1552 => x"9386f6ff",
        1553 => x"3377d700",
        1554 => x"13170701",
        1555 => x"b3fede00",
        1556 => x"3307d701",
        1557 => x"63e6f500",
        1558 => x"639ef500",
        1559 => x"637ce500",
        1560 => x"3306c740",
        1561 => x"3337c700",
        1562 => x"33076700",
        1563 => x"b387e740",
        1564 => x"13070600",
        1565 => x"3307e540",
        1566 => x"3335e500",
        1567 => x"b385f540",
        1568 => x"b385a540",
        1569 => x"b3981501",
        1570 => x"33570701",
        1571 => x"33e5e800",
        1572 => x"b3d50501",
        1573 => x"67800000",
        1574 => x"13030500",
        1575 => x"630e0600",
        1576 => x"83830500",
        1577 => x"23007300",
        1578 => x"1306f6ff",
        1579 => x"13031300",
        1580 => x"93851500",
        1581 => x"e31606fe",
        1582 => x"67800000",
        1583 => x"13030500",
        1584 => x"630a0600",
        1585 => x"2300b300",
        1586 => x"1306f6ff",
        1587 => x"13031300",
        1588 => x"e31a06fe",
        1589 => x"67800000",
        1590 => x"630c0602",
        1591 => x"13030500",
        1592 => x"93061000",
        1593 => x"636ab500",
        1594 => x"9306f0ff",
        1595 => x"1307f6ff",
        1596 => x"3303e300",
        1597 => x"b385e500",
        1598 => x"83830500",
        1599 => x"23007300",
        1600 => x"1306f6ff",
        1601 => x"3303d300",
        1602 => x"b385d500",
        1603 => x"e31606fe",
        1604 => x"67800000",
        1605 => x"130101f9",
        1606 => x"23248106",
        1607 => x"232e3105",
        1608 => x"23261106",
        1609 => x"23229106",
        1610 => x"23202107",
        1611 => x"232c4105",
        1612 => x"232a5105",
        1613 => x"23286105",
        1614 => x"23267105",
        1615 => x"23248105",
        1616 => x"93090500",
        1617 => x"13840500",
        1618 => x"232c0100",
        1619 => x"232e0100",
        1620 => x"23200102",
        1621 => x"23220102",
        1622 => x"23240102",
        1623 => x"23260102",
        1624 => x"23280102",
        1625 => x"232a0102",
        1626 => x"232c0102",
        1627 => x"232e0102",
        1628 => x"97f2ffff",
        1629 => x"93821296",
        1630 => x"73905230",
        1631 => x"b7220000",
        1632 => x"93828280",
        1633 => x"73900230",
        1634 => x"efe04fef",
        1635 => x"b7877d01",
        1636 => x"370700f0",
        1637 => x"9387f783",
        1638 => x"2326f708",
        1639 => x"37390000",
        1640 => x"93071001",
        1641 => x"2320f708",
        1642 => x"13054920",
        1643 => x"efe08ff0",
        1644 => x"63543003",
        1645 => x"9384f9ff",
        1646 => x"9309f0ff",
        1647 => x"03250400",
        1648 => x"9384f4ff",
        1649 => x"13044400",
        1650 => x"efe0cfee",
        1651 => x"13054920",
        1652 => x"efe04fee",
        1653 => x"e39434ff",
        1654 => x"37350000",
        1655 => x"1305851d",
        1656 => x"371a0000",
        1657 => x"b71b0000",
        1658 => x"efe0cfec",
        1659 => x"13040000",
        1660 => x"373c0000",
        1661 => x"130a0ae1",
        1662 => x"930a0000",
        1663 => x"938b0bfa",
        1664 => x"93050000",
        1665 => x"13058100",
        1666 => x"ef00c026",
        1667 => x"13041400",
        1668 => x"63020502",
        1669 => x"e31674ff",
        1670 => x"73001000",
        1671 => x"93050000",
        1672 => x"13058100",
        1673 => x"13040000",
        1674 => x"ef00c024",
        1675 => x"13041400",
        1676 => x"e31205fe",
        1677 => x"83248100",
        1678 => x"032bc100",
        1679 => x"1306c003",
        1680 => x"93060000",
        1681 => x"13850400",
        1682 => x"93050b00",
        1683 => x"eff08f9e",
        1684 => x"93090500",
        1685 => x"1306c003",
        1686 => x"93060000",
        1687 => x"13850400",
        1688 => x"93050b00",
        1689 => x"efe09fd5",
        1690 => x"1306c003",
        1691 => x"93060000",
        1692 => x"eff04f9c",
        1693 => x"13060a00",
        1694 => x"93860a00",
        1695 => x"13090500",
        1696 => x"93050b00",
        1697 => x"13850400",
        1698 => x"efe05fd3",
        1699 => x"83260101",
        1700 => x"13070500",
        1701 => x"13880900",
        1702 => x"93070900",
        1703 => x"13860400",
        1704 => x"93058c20",
        1705 => x"13058101",
        1706 => x"ef00c015",
        1707 => x"13058101",
        1708 => x"efe04fe0",
        1709 => x"e31674f5",
        1710 => x"6ff01ff6",
        1711 => x"03a5c187",
        1712 => x"67800000",
        1713 => x"130101ff",
        1714 => x"23248100",
        1715 => x"23261100",
        1716 => x"93070000",
        1717 => x"13040500",
        1718 => x"63880700",
        1719 => x"93050000",
        1720 => x"97000000",
        1721 => x"e7000000",
        1722 => x"b7370000",
        1723 => x"03a58737",
        1724 => x"83278502",
        1725 => x"63840700",
        1726 => x"e7800700",
        1727 => x"13050400",
        1728 => x"ef108033",
        1729 => x"130101ff",
        1730 => x"23248100",
        1731 => x"23229100",
        1732 => x"37340000",
        1733 => x"b7340000",
        1734 => x"9387c437",
        1735 => x"1304c437",
        1736 => x"3304f440",
        1737 => x"23202101",
        1738 => x"23261100",
        1739 => x"13542440",
        1740 => x"9384c437",
        1741 => x"13090000",
        1742 => x"63108904",
        1743 => x"b7340000",
        1744 => x"37340000",
        1745 => x"9387c437",
        1746 => x"1304c437",
        1747 => x"3304f440",
        1748 => x"13542440",
        1749 => x"9384c437",
        1750 => x"13090000",
        1751 => x"63188902",
        1752 => x"8320c100",
        1753 => x"03248100",
        1754 => x"83244100",
        1755 => x"03290100",
        1756 => x"13010101",
        1757 => x"67800000",
        1758 => x"83a70400",
        1759 => x"13091900",
        1760 => x"93844400",
        1761 => x"e7800700",
        1762 => x"6ff01ffb",
        1763 => x"83a70400",
        1764 => x"13091900",
        1765 => x"93844400",
        1766 => x"e7800700",
        1767 => x"6ff01ffc",
        1768 => x"130101f6",
        1769 => x"232af108",
        1770 => x"b7070080",
        1771 => x"93c7f7ff",
        1772 => x"232ef100",
        1773 => x"2328f100",
        1774 => x"b707ffff",
        1775 => x"2326d108",
        1776 => x"2324b100",
        1777 => x"232cb100",
        1778 => x"93878720",
        1779 => x"9306c108",
        1780 => x"93058100",
        1781 => x"232e1106",
        1782 => x"232af100",
        1783 => x"2328e108",
        1784 => x"232c0109",
        1785 => x"232e1109",
        1786 => x"2322d100",
        1787 => x"ef004041",
        1788 => x"83278100",
        1789 => x"23800700",
        1790 => x"8320c107",
        1791 => x"1301010a",
        1792 => x"67800000",
        1793 => x"130101f6",
        1794 => x"232af108",
        1795 => x"b7070080",
        1796 => x"93c7f7ff",
        1797 => x"232ef100",
        1798 => x"2328f100",
        1799 => x"b707ffff",
        1800 => x"93878720",
        1801 => x"232af100",
        1802 => x"2324a100",
        1803 => x"232ca100",
        1804 => x"03a5c187",
        1805 => x"2324c108",
        1806 => x"2326d108",
        1807 => x"13860500",
        1808 => x"93068108",
        1809 => x"93058100",
        1810 => x"232e1106",
        1811 => x"2328e108",
        1812 => x"232c0109",
        1813 => x"232e1109",
        1814 => x"2322d100",
        1815 => x"ef00403a",
        1816 => x"83278100",
        1817 => x"23800700",
        1818 => x"8320c107",
        1819 => x"1301010a",
        1820 => x"67800000",
        1821 => x"13860500",
        1822 => x"93050500",
        1823 => x"03a5c187",
        1824 => x"6f004000",
        1825 => x"130101ff",
        1826 => x"23248100",
        1827 => x"23229100",
        1828 => x"13040500",
        1829 => x"13850500",
        1830 => x"93050600",
        1831 => x"23261100",
        1832 => x"23a20188",
        1833 => x"ef10401c",
        1834 => x"9307f0ff",
        1835 => x"6318f500",
        1836 => x"83a74188",
        1837 => x"63840700",
        1838 => x"2320f400",
        1839 => x"8320c100",
        1840 => x"03248100",
        1841 => x"83244100",
        1842 => x"13010101",
        1843 => x"67800000",
        1844 => x"130101fe",
        1845 => x"23282101",
        1846 => x"03a98500",
        1847 => x"232c8100",
        1848 => x"23263101",
        1849 => x"23244101",
        1850 => x"23225101",
        1851 => x"232e1100",
        1852 => x"232a9100",
        1853 => x"23206101",
        1854 => x"83aa0500",
        1855 => x"13840500",
        1856 => x"130a0600",
        1857 => x"93890600",
        1858 => x"63ec2609",
        1859 => x"83d7c500",
        1860 => x"13f70748",
        1861 => x"63040708",
        1862 => x"03274401",
        1863 => x"93043000",
        1864 => x"83a50501",
        1865 => x"b384e402",
        1866 => x"13072000",
        1867 => x"b38aba40",
        1868 => x"130b0500",
        1869 => x"b3c4e402",
        1870 => x"13871600",
        1871 => x"33075701",
        1872 => x"63f4e400",
        1873 => x"93040700",
        1874 => x"93f70740",
        1875 => x"6386070a",
        1876 => x"93850400",
        1877 => x"13050b00",
        1878 => x"ef001065",
        1879 => x"13090500",
        1880 => x"630c050a",
        1881 => x"83250401",
        1882 => x"13860a00",
        1883 => x"eff0dfb2",
        1884 => x"8357c400",
        1885 => x"93f7f7b7",
        1886 => x"93e70708",
        1887 => x"2316f400",
        1888 => x"23282401",
        1889 => x"232a9400",
        1890 => x"33095901",
        1891 => x"b3845441",
        1892 => x"23202401",
        1893 => x"23249400",
        1894 => x"13890900",
        1895 => x"63f42901",
        1896 => x"13890900",
        1897 => x"03250400",
        1898 => x"13060900",
        1899 => x"93050a00",
        1900 => x"eff09fb2",
        1901 => x"83278400",
        1902 => x"13050000",
        1903 => x"b3872741",
        1904 => x"2324f400",
        1905 => x"83270400",
        1906 => x"b3872701",
        1907 => x"2320f400",
        1908 => x"8320c101",
        1909 => x"03248101",
        1910 => x"83244101",
        1911 => x"03290101",
        1912 => x"8329c100",
        1913 => x"032a8100",
        1914 => x"832a4100",
        1915 => x"032b0100",
        1916 => x"13010102",
        1917 => x"67800000",
        1918 => x"13860400",
        1919 => x"13050b00",
        1920 => x"ef00906f",
        1921 => x"13090500",
        1922 => x"e31c05f6",
        1923 => x"83250401",
        1924 => x"13050b00",
        1925 => x"ef00d049",
        1926 => x"9307c000",
        1927 => x"2320fb00",
        1928 => x"8357c400",
        1929 => x"1305f0ff",
        1930 => x"93e70704",
        1931 => x"2316f400",
        1932 => x"6ff01ffa",
        1933 => x"83278600",
        1934 => x"130101fd",
        1935 => x"232e3101",
        1936 => x"23286101",
        1937 => x"23261102",
        1938 => x"23248102",
        1939 => x"23229102",
        1940 => x"23202103",
        1941 => x"232c4101",
        1942 => x"232a5101",
        1943 => x"23267101",
        1944 => x"23248101",
        1945 => x"23229101",
        1946 => x"2320a101",
        1947 => x"032b0600",
        1948 => x"93090600",
        1949 => x"63980712",
        1950 => x"13050000",
        1951 => x"8320c102",
        1952 => x"03248102",
        1953 => x"23a20900",
        1954 => x"83244102",
        1955 => x"03290102",
        1956 => x"8329c101",
        1957 => x"032a8101",
        1958 => x"832a4101",
        1959 => x"032b0101",
        1960 => x"832bc100",
        1961 => x"032c8100",
        1962 => x"832c4100",
        1963 => x"032d0100",
        1964 => x"13010103",
        1965 => x"67800000",
        1966 => x"832a0b00",
        1967 => x"032d4b00",
        1968 => x"130b8b00",
        1969 => x"03298400",
        1970 => x"832c0400",
        1971 => x"e3060dfe",
        1972 => x"63642d09",
        1973 => x"8357c400",
        1974 => x"13f70748",
        1975 => x"630e0706",
        1976 => x"83244401",
        1977 => x"83250401",
        1978 => x"b3849b02",
        1979 => x"b38cbc40",
        1980 => x"13871c00",
        1981 => x"3307a701",
        1982 => x"b3c48403",
        1983 => x"63f4e400",
        1984 => x"93040700",
        1985 => x"93f70740",
        1986 => x"638c070a",
        1987 => x"93850400",
        1988 => x"13050a00",
        1989 => x"ef005049",
        1990 => x"13090500",
        1991 => x"6302050c",
        1992 => x"83250401",
        1993 => x"13860c00",
        1994 => x"eff01f97",
        1995 => x"8357c400",
        1996 => x"93f7f7b7",
        1997 => x"93e70708",
        1998 => x"2316f400",
        1999 => x"23282401",
        2000 => x"232a9400",
        2001 => x"33099901",
        2002 => x"b3849441",
        2003 => x"23202401",
        2004 => x"23249400",
        2005 => x"13090d00",
        2006 => x"63742d01",
        2007 => x"13090d00",
        2008 => x"03250400",
        2009 => x"93850a00",
        2010 => x"13060900",
        2011 => x"eff0df96",
        2012 => x"83278400",
        2013 => x"b38aaa01",
        2014 => x"b3872741",
        2015 => x"2324f400",
        2016 => x"83270400",
        2017 => x"b3872701",
        2018 => x"2320f400",
        2019 => x"83a78900",
        2020 => x"b387a741",
        2021 => x"23a4f900",
        2022 => x"e38007ee",
        2023 => x"130d0000",
        2024 => x"6ff05ff2",
        2025 => x"130a0500",
        2026 => x"13840500",
        2027 => x"930a0000",
        2028 => x"130d0000",
        2029 => x"930b3000",
        2030 => x"130c2000",
        2031 => x"6ff09ff0",
        2032 => x"13860400",
        2033 => x"13050a00",
        2034 => x"ef001053",
        2035 => x"13090500",
        2036 => x"e31605f6",
        2037 => x"83250401",
        2038 => x"13050a00",
        2039 => x"ef00502d",
        2040 => x"9307c000",
        2041 => x"2320fa00",
        2042 => x"8357c400",
        2043 => x"1305f0ff",
        2044 => x"93e70704",
        2045 => x"2316f400",
        2046 => x"23a40900",
        2047 => x"6ff01fe8",
        2048 => x"83d7c500",
        2049 => x"130101f5",
        2050 => x"2324810a",
        2051 => x"2322910a",
        2052 => x"2320210b",
        2053 => x"232c4109",
        2054 => x"2326110a",
        2055 => x"232e3109",
        2056 => x"232a5109",
        2057 => x"23286109",
        2058 => x"23267109",
        2059 => x"23248109",
        2060 => x"23229109",
        2061 => x"2320a109",
        2062 => x"232eb107",
        2063 => x"93f70708",
        2064 => x"130a0500",
        2065 => x"13890500",
        2066 => x"93040600",
        2067 => x"13840600",
        2068 => x"63880706",
        2069 => x"83a70501",
        2070 => x"63940706",
        2071 => x"93050004",
        2072 => x"ef009034",
        2073 => x"2320a900",
        2074 => x"2328a900",
        2075 => x"63160504",
        2076 => x"9307c000",
        2077 => x"2320fa00",
        2078 => x"1305f0ff",
        2079 => x"8320c10a",
        2080 => x"0324810a",
        2081 => x"8324410a",
        2082 => x"0329010a",
        2083 => x"8329c109",
        2084 => x"032a8109",
        2085 => x"832a4109",
        2086 => x"032b0109",
        2087 => x"832bc108",
        2088 => x"032c8108",
        2089 => x"832c4108",
        2090 => x"032d0108",
        2091 => x"832dc107",
        2092 => x"1301010b",
        2093 => x"67800000",
        2094 => x"93070004",
        2095 => x"232af900",
        2096 => x"93070002",
        2097 => x"a304f102",
        2098 => x"93070003",
        2099 => x"23220102",
        2100 => x"2305f102",
        2101 => x"23268100",
        2102 => x"930c5002",
        2103 => x"373b0000",
        2104 => x"b73b0000",
        2105 => x"373d0000",
        2106 => x"372c0000",
        2107 => x"930a0000",
        2108 => x"13840400",
        2109 => x"83470400",
        2110 => x"63840700",
        2111 => x"639c970d",
        2112 => x"b30d9440",
        2113 => x"63069402",
        2114 => x"93860d00",
        2115 => x"13860400",
        2116 => x"93050900",
        2117 => x"13050a00",
        2118 => x"eff09fbb",
        2119 => x"9307f0ff",
        2120 => x"6306f524",
        2121 => x"83274102",
        2122 => x"b387b701",
        2123 => x"2322f102",
        2124 => x"83470400",
        2125 => x"638c0722",
        2126 => x"9307f0ff",
        2127 => x"93041400",
        2128 => x"23280100",
        2129 => x"232e0100",
        2130 => x"232af100",
        2131 => x"232c0100",
        2132 => x"a3090104",
        2133 => x"23240106",
        2134 => x"930d1000",
        2135 => x"83c50400",
        2136 => x"13065000",
        2137 => x"13054b2e",
        2138 => x"ef005012",
        2139 => x"83270101",
        2140 => x"13841400",
        2141 => x"63140506",
        2142 => x"13f70701",
        2143 => x"63060700",
        2144 => x"13070002",
        2145 => x"a309e104",
        2146 => x"13f78700",
        2147 => x"63060700",
        2148 => x"1307b002",
        2149 => x"a309e104",
        2150 => x"83c60400",
        2151 => x"1307a002",
        2152 => x"638ce604",
        2153 => x"8327c101",
        2154 => x"13840400",
        2155 => x"93060000",
        2156 => x"13069000",
        2157 => x"1305a000",
        2158 => x"03470400",
        2159 => x"93051400",
        2160 => x"130707fd",
        2161 => x"637ce608",
        2162 => x"63840604",
        2163 => x"232ef100",
        2164 => x"6f000004",
        2165 => x"13041400",
        2166 => x"6ff0dff1",
        2167 => x"13074b2e",
        2168 => x"3305e540",
        2169 => x"3395ad00",
        2170 => x"b3e7a700",
        2171 => x"2328f100",
        2172 => x"93040400",
        2173 => x"6ff09ff6",
        2174 => x"0327c100",
        2175 => x"93064700",
        2176 => x"03270700",
        2177 => x"2326d100",
        2178 => x"63400704",
        2179 => x"232ee100",
        2180 => x"03470400",
        2181 => x"9307e002",
        2182 => x"6316f708",
        2183 => x"03471400",
        2184 => x"9307a002",
        2185 => x"631af704",
        2186 => x"8327c100",
        2187 => x"13042400",
        2188 => x"13874700",
        2189 => x"83a70700",
        2190 => x"2326e100",
        2191 => x"63ca0702",
        2192 => x"232af100",
        2193 => x"6f000006",
        2194 => x"3307e040",
        2195 => x"93e72700",
        2196 => x"232ee100",
        2197 => x"2328f100",
        2198 => x"6ff09ffb",
        2199 => x"b387a702",
        2200 => x"13840500",
        2201 => x"93061000",
        2202 => x"b387e700",
        2203 => x"6ff0dff4",
        2204 => x"9307f0ff",
        2205 => x"6ff0dffc",
        2206 => x"13041400",
        2207 => x"232a0100",
        2208 => x"93060000",
        2209 => x"93070000",
        2210 => x"13069000",
        2211 => x"1305a000",
        2212 => x"03470400",
        2213 => x"93051400",
        2214 => x"130707fd",
        2215 => x"6372e608",
        2216 => x"e39006fa",
        2217 => x"83450400",
        2218 => x"13063000",
        2219 => x"1385cb2e",
        2220 => x"ef00c07d",
        2221 => x"63020502",
        2222 => x"9387cb2e",
        2223 => x"3305f540",
        2224 => x"83270101",
        2225 => x"13070004",
        2226 => x"3317a700",
        2227 => x"b3e7e700",
        2228 => x"13041400",
        2229 => x"2328f100",
        2230 => x"83450400",
        2231 => x"13066000",
        2232 => x"13050d2f",
        2233 => x"93041400",
        2234 => x"2304b102",
        2235 => x"ef00007a",
        2236 => x"630a0508",
        2237 => x"63980a04",
        2238 => x"03270101",
        2239 => x"8327c100",
        2240 => x"13770710",
        2241 => x"63080702",
        2242 => x"93874700",
        2243 => x"2326f100",
        2244 => x"83274102",
        2245 => x"b3873701",
        2246 => x"2322f102",
        2247 => x"6ff05fdd",
        2248 => x"b387a702",
        2249 => x"13840500",
        2250 => x"93061000",
        2251 => x"b387e700",
        2252 => x"6ff01ff6",
        2253 => x"93877700",
        2254 => x"93f787ff",
        2255 => x"93878700",
        2256 => x"6ff0dffc",
        2257 => x"1307c100",
        2258 => x"93060ccd",
        2259 => x"13060900",
        2260 => x"93050101",
        2261 => x"13050a00",
        2262 => x"97000000",
        2263 => x"e7000000",
        2264 => x"9307f0ff",
        2265 => x"93090500",
        2266 => x"e314f5fa",
        2267 => x"8357c900",
        2268 => x"1305f0ff",
        2269 => x"93f70704",
        2270 => x"e39207d0",
        2271 => x"03254102",
        2272 => x"6ff0dfcf",
        2273 => x"1307c100",
        2274 => x"93060ccd",
        2275 => x"13060900",
        2276 => x"93050101",
        2277 => x"13050a00",
        2278 => x"ef00801b",
        2279 => x"6ff05ffc",
        2280 => x"130101fd",
        2281 => x"232c4101",
        2282 => x"83a70501",
        2283 => x"130a0700",
        2284 => x"03a78500",
        2285 => x"23248102",
        2286 => x"23202103",
        2287 => x"232e3101",
        2288 => x"232a5101",
        2289 => x"23261102",
        2290 => x"23229102",
        2291 => x"23286101",
        2292 => x"23267101",
        2293 => x"93090500",
        2294 => x"13840500",
        2295 => x"13090600",
        2296 => x"938a0600",
        2297 => x"63d4e700",
        2298 => x"93070700",
        2299 => x"2320f900",
        2300 => x"03473404",
        2301 => x"63060700",
        2302 => x"93871700",
        2303 => x"2320f900",
        2304 => x"83270400",
        2305 => x"93f70702",
        2306 => x"63880700",
        2307 => x"83270900",
        2308 => x"93872700",
        2309 => x"2320f900",
        2310 => x"83240400",
        2311 => x"93f46400",
        2312 => x"639e0400",
        2313 => x"130b9401",
        2314 => x"930bf0ff",
        2315 => x"8327c400",
        2316 => x"03270900",
        2317 => x"b387e740",
        2318 => x"63c2f408",
        2319 => x"83473404",
        2320 => x"b336f000",
        2321 => x"83270400",
        2322 => x"93f70702",
        2323 => x"6390070c",
        2324 => x"13063404",
        2325 => x"93850a00",
        2326 => x"13850900",
        2327 => x"e7000a00",
        2328 => x"9307f0ff",
        2329 => x"6308f506",
        2330 => x"83270400",
        2331 => x"13074000",
        2332 => x"93040000",
        2333 => x"93f76700",
        2334 => x"639ce700",
        2335 => x"8324c400",
        2336 => x"83270900",
        2337 => x"b384f440",
        2338 => x"63d40400",
        2339 => x"93040000",
        2340 => x"83278400",
        2341 => x"03270401",
        2342 => x"6356f700",
        2343 => x"b387e740",
        2344 => x"b384f400",
        2345 => x"13090000",
        2346 => x"1304a401",
        2347 => x"130bf0ff",
        2348 => x"63902409",
        2349 => x"13050000",
        2350 => x"6f000002",
        2351 => x"93061000",
        2352 => x"13060b00",
        2353 => x"93850a00",
        2354 => x"13850900",
        2355 => x"e7000a00",
        2356 => x"631a7503",
        2357 => x"1305f0ff",
        2358 => x"8320c102",
        2359 => x"03248102",
        2360 => x"83244102",
        2361 => x"03290102",
        2362 => x"8329c101",
        2363 => x"032a8101",
        2364 => x"832a4101",
        2365 => x"032b0101",
        2366 => x"832bc100",
        2367 => x"13010103",
        2368 => x"67800000",
        2369 => x"93841400",
        2370 => x"6ff05ff2",
        2371 => x"3307d400",
        2372 => x"13060003",
        2373 => x"a301c704",
        2374 => x"03475404",
        2375 => x"93871600",
        2376 => x"b307f400",
        2377 => x"93862600",
        2378 => x"a381e704",
        2379 => x"6ff05ff2",
        2380 => x"93061000",
        2381 => x"13060400",
        2382 => x"93850a00",
        2383 => x"13850900",
        2384 => x"e7000a00",
        2385 => x"e30865f9",
        2386 => x"13091900",
        2387 => x"6ff05ff6",
        2388 => x"130101fd",
        2389 => x"23248102",
        2390 => x"23229102",
        2391 => x"23202103",
        2392 => x"232e3101",
        2393 => x"23261102",
        2394 => x"232c4101",
        2395 => x"232a5101",
        2396 => x"23286101",
        2397 => x"83c88501",
        2398 => x"93078007",
        2399 => x"93040500",
        2400 => x"13840500",
        2401 => x"13090600",
        2402 => x"93890600",
        2403 => x"63ee1701",
        2404 => x"93072006",
        2405 => x"93863504",
        2406 => x"63ee1701",
        2407 => x"63840828",
        2408 => x"93078005",
        2409 => x"6388f822",
        2410 => x"930a2404",
        2411 => x"23011405",
        2412 => x"6f004004",
        2413 => x"9387d8f9",
        2414 => x"93f7f70f",
        2415 => x"13065001",
        2416 => x"e364f6fe",
        2417 => x"37360000",
        2418 => x"93972700",
        2419 => x"13060632",
        2420 => x"b387c700",
        2421 => x"83a70700",
        2422 => x"67800700",
        2423 => x"83270700",
        2424 => x"938a2504",
        2425 => x"93864700",
        2426 => x"83a70700",
        2427 => x"2320d700",
        2428 => x"2381f504",
        2429 => x"93071000",
        2430 => x"6f008026",
        2431 => x"83a70500",
        2432 => x"03250700",
        2433 => x"13f60708",
        2434 => x"93054500",
        2435 => x"63060602",
        2436 => x"83270500",
        2437 => x"2320b700",
        2438 => x"37380000",
        2439 => x"63d80700",
        2440 => x"1307d002",
        2441 => x"b307f040",
        2442 => x"a301e404",
        2443 => x"1308882f",
        2444 => x"1307a000",
        2445 => x"6f008006",
        2446 => x"13f60704",
        2447 => x"83270500",
        2448 => x"2320b700",
        2449 => x"e30a06fc",
        2450 => x"93970701",
        2451 => x"93d70741",
        2452 => x"6ff09ffc",
        2453 => x"03a60500",
        2454 => x"83270700",
        2455 => x"13750608",
        2456 => x"93854700",
        2457 => x"63080500",
        2458 => x"2320b700",
        2459 => x"83a70700",
        2460 => x"6f004001",
        2461 => x"13760604",
        2462 => x"2320b700",
        2463 => x"e30806fe",
        2464 => x"83d70700",
        2465 => x"37380000",
        2466 => x"1307f006",
        2467 => x"1308882f",
        2468 => x"6388e814",
        2469 => x"1307a000",
        2470 => x"a3010404",
        2471 => x"03264400",
        2472 => x"2324c400",
        2473 => x"63480600",
        2474 => x"83250400",
        2475 => x"93f5b5ff",
        2476 => x"2320b400",
        2477 => x"63960700",
        2478 => x"938a0600",
        2479 => x"63040602",
        2480 => x"938a0600",
        2481 => x"33f6e702",
        2482 => x"938afaff",
        2483 => x"3306c800",
        2484 => x"03460600",
        2485 => x"2380ca00",
        2486 => x"13860700",
        2487 => x"b3d7e702",
        2488 => x"e372e6fe",
        2489 => x"93078000",
        2490 => x"6314f702",
        2491 => x"83270400",
        2492 => x"93f71700",
        2493 => x"638e0700",
        2494 => x"03274400",
        2495 => x"83270401",
        2496 => x"63c8e700",
        2497 => x"93070003",
        2498 => x"a38ffafe",
        2499 => x"938afaff",
        2500 => x"b3865641",
        2501 => x"2328d400",
        2502 => x"13870900",
        2503 => x"93060900",
        2504 => x"1306c100",
        2505 => x"93050400",
        2506 => x"13850400",
        2507 => x"eff05fc7",
        2508 => x"130af0ff",
        2509 => x"631c4513",
        2510 => x"1305f0ff",
        2511 => x"8320c102",
        2512 => x"03248102",
        2513 => x"83244102",
        2514 => x"03290102",
        2515 => x"8329c101",
        2516 => x"032a8101",
        2517 => x"832a4101",
        2518 => x"032b0101",
        2519 => x"13010103",
        2520 => x"67800000",
        2521 => x"83a70500",
        2522 => x"93e70702",
        2523 => x"23a0f500",
        2524 => x"37380000",
        2525 => x"93088007",
        2526 => x"1308c830",
        2527 => x"a3021405",
        2528 => x"03260400",
        2529 => x"83250700",
        2530 => x"13750608",
        2531 => x"83a70500",
        2532 => x"93854500",
        2533 => x"631a0500",
        2534 => x"13750604",
        2535 => x"63060500",
        2536 => x"93970701",
        2537 => x"93d70701",
        2538 => x"2320b700",
        2539 => x"13771600",
        2540 => x"63060700",
        2541 => x"13660602",
        2542 => x"2320c400",
        2543 => x"13070001",
        2544 => x"e39c07ec",
        2545 => x"03260400",
        2546 => x"1376f6fd",
        2547 => x"2320c400",
        2548 => x"6ff09fec",
        2549 => x"37380000",
        2550 => x"1308882f",
        2551 => x"6ff01ffa",
        2552 => x"13078000",
        2553 => x"6ff05feb",
        2554 => x"03a60500",
        2555 => x"83270700",
        2556 => x"83a54501",
        2557 => x"13780608",
        2558 => x"13854700",
        2559 => x"630a0800",
        2560 => x"2320a700",
        2561 => x"83a70700",
        2562 => x"23a0b700",
        2563 => x"6f008001",
        2564 => x"2320a700",
        2565 => x"13760604",
        2566 => x"83a70700",
        2567 => x"e30606fe",
        2568 => x"2390b700",
        2569 => x"23280400",
        2570 => x"938a0600",
        2571 => x"6ff0dfee",
        2572 => x"83270700",
        2573 => x"03a64500",
        2574 => x"93050000",
        2575 => x"93864700",
        2576 => x"2320d700",
        2577 => x"83aa0700",
        2578 => x"13850a00",
        2579 => x"ef000024",
        2580 => x"63060500",
        2581 => x"33055541",
        2582 => x"2322a400",
        2583 => x"83274400",
        2584 => x"2328f400",
        2585 => x"a3010404",
        2586 => x"6ff01feb",
        2587 => x"83260401",
        2588 => x"13860a00",
        2589 => x"93050900",
        2590 => x"13850400",
        2591 => x"e7800900",
        2592 => x"e30c45eb",
        2593 => x"83270400",
        2594 => x"93f72700",
        2595 => x"63940704",
        2596 => x"8327c100",
        2597 => x"0325c400",
        2598 => x"e352f5ea",
        2599 => x"13850700",
        2600 => x"6ff0dfe9",
        2601 => x"93061000",
        2602 => x"13860a00",
        2603 => x"93050900",
        2604 => x"13850400",
        2605 => x"e7800900",
        2606 => x"e30065e9",
        2607 => x"130a1a00",
        2608 => x"8327c400",
        2609 => x"0327c100",
        2610 => x"b387e740",
        2611 => x"e34cfafc",
        2612 => x"6ff01ffc",
        2613 => x"130a0000",
        2614 => x"930a9401",
        2615 => x"130bf0ff",
        2616 => x"6ff01ffe",
        2617 => x"130101ff",
        2618 => x"23248100",
        2619 => x"13840500",
        2620 => x"83a50500",
        2621 => x"23229100",
        2622 => x"23261100",
        2623 => x"93040500",
        2624 => x"63840500",
        2625 => x"eff01ffe",
        2626 => x"93050400",
        2627 => x"03248100",
        2628 => x"8320c100",
        2629 => x"13850400",
        2630 => x"83244100",
        2631 => x"13010101",
        2632 => x"6f000019",
        2633 => x"83a7c187",
        2634 => x"6380a716",
        2635 => x"83274502",
        2636 => x"130101fe",
        2637 => x"232c8100",
        2638 => x"232e1100",
        2639 => x"232a9100",
        2640 => x"23282101",
        2641 => x"23263101",
        2642 => x"13040500",
        2643 => x"63840702",
        2644 => x"83a7c700",
        2645 => x"93040000",
        2646 => x"13090008",
        2647 => x"6392070e",
        2648 => x"83274402",
        2649 => x"83a50700",
        2650 => x"63860500",
        2651 => x"13050400",
        2652 => x"ef000014",
        2653 => x"83254401",
        2654 => x"63860500",
        2655 => x"13050400",
        2656 => x"ef000013",
        2657 => x"83254402",
        2658 => x"63860500",
        2659 => x"13050400",
        2660 => x"ef000012",
        2661 => x"83258403",
        2662 => x"63860500",
        2663 => x"13050400",
        2664 => x"ef000011",
        2665 => x"8325c403",
        2666 => x"63860500",
        2667 => x"13050400",
        2668 => x"ef000010",
        2669 => x"83250404",
        2670 => x"63860500",
        2671 => x"13050400",
        2672 => x"ef00000f",
        2673 => x"8325c405",
        2674 => x"63860500",
        2675 => x"13050400",
        2676 => x"ef00000e",
        2677 => x"83258405",
        2678 => x"63860500",
        2679 => x"13050400",
        2680 => x"ef00000d",
        2681 => x"83254403",
        2682 => x"63860500",
        2683 => x"13050400",
        2684 => x"ef00000c",
        2685 => x"83278401",
        2686 => x"638a0706",
        2687 => x"83278402",
        2688 => x"13050400",
        2689 => x"e7800700",
        2690 => x"83258404",
        2691 => x"63800506",
        2692 => x"13050400",
        2693 => x"03248101",
        2694 => x"8320c101",
        2695 => x"83244101",
        2696 => x"03290101",
        2697 => x"8329c100",
        2698 => x"13010102",
        2699 => x"6ff09feb",
        2700 => x"b3859500",
        2701 => x"83a50500",
        2702 => x"63900502",
        2703 => x"93844400",
        2704 => x"83274402",
        2705 => x"83a5c700",
        2706 => x"e39424ff",
        2707 => x"13050400",
        2708 => x"ef000006",
        2709 => x"6ff0dff0",
        2710 => x"83a90500",
        2711 => x"13050400",
        2712 => x"ef000005",
        2713 => x"93850900",
        2714 => x"6ff01ffd",
        2715 => x"8320c101",
        2716 => x"03248101",
        2717 => x"83244101",
        2718 => x"03290101",
        2719 => x"8329c100",
        2720 => x"13010102",
        2721 => x"67800000",
        2722 => x"67800000",
        2723 => x"93f5f50f",
        2724 => x"3306c500",
        2725 => x"6316c500",
        2726 => x"13050000",
        2727 => x"67800000",
        2728 => x"83470500",
        2729 => x"e38cb7fe",
        2730 => x"13051500",
        2731 => x"6ff09ffe",
        2732 => x"638a050e",
        2733 => x"83a7c5ff",
        2734 => x"130101fe",
        2735 => x"232c8100",
        2736 => x"232e1100",
        2737 => x"1384c5ff",
        2738 => x"63d40700",
        2739 => x"3304f400",
        2740 => x"2326a100",
        2741 => x"ef000034",
        2742 => x"83a78188",
        2743 => x"0325c100",
        2744 => x"639e0700",
        2745 => x"23220400",
        2746 => x"23a48188",
        2747 => x"03248101",
        2748 => x"8320c101",
        2749 => x"13010102",
        2750 => x"6f000032",
        2751 => x"6374f402",
        2752 => x"03260400",
        2753 => x"b306c400",
        2754 => x"639ad700",
        2755 => x"83a60700",
        2756 => x"83a74700",
        2757 => x"b386c600",
        2758 => x"2320d400",
        2759 => x"2322f400",
        2760 => x"6ff09ffc",
        2761 => x"13870700",
        2762 => x"83a74700",
        2763 => x"63840700",
        2764 => x"e37af4fe",
        2765 => x"83260700",
        2766 => x"3306d700",
        2767 => x"63188602",
        2768 => x"03260400",
        2769 => x"b386c600",
        2770 => x"2320d700",
        2771 => x"3306d700",
        2772 => x"e39ec7f8",
        2773 => x"03a60700",
        2774 => x"83a74700",
        2775 => x"b306d600",
        2776 => x"2320d700",
        2777 => x"2322f700",
        2778 => x"6ff05ff8",
        2779 => x"6378c400",
        2780 => x"9307c000",
        2781 => x"2320f500",
        2782 => x"6ff05ff7",
        2783 => x"03260400",
        2784 => x"b306c400",
        2785 => x"639ad700",
        2786 => x"83a60700",
        2787 => x"83a74700",
        2788 => x"b386c600",
        2789 => x"2320d400",
        2790 => x"2322f400",
        2791 => x"23228700",
        2792 => x"6ff0dff4",
        2793 => x"67800000",
        2794 => x"130101fe",
        2795 => x"232a9100",
        2796 => x"93843500",
        2797 => x"93f4c4ff",
        2798 => x"23282101",
        2799 => x"232e1100",
        2800 => x"232c8100",
        2801 => x"23263101",
        2802 => x"93848400",
        2803 => x"9307c000",
        2804 => x"13090500",
        2805 => x"63f4f406",
        2806 => x"9304c000",
        2807 => x"63e2b406",
        2808 => x"13050900",
        2809 => x"ef000023",
        2810 => x"03a78188",
        2811 => x"93868188",
        2812 => x"13040700",
        2813 => x"631a0406",
        2814 => x"1384c188",
        2815 => x"83270400",
        2816 => x"639a0700",
        2817 => x"93050000",
        2818 => x"13050900",
        2819 => x"ef00001c",
        2820 => x"2320a400",
        2821 => x"93850400",
        2822 => x"13050900",
        2823 => x"ef00001b",
        2824 => x"9309f0ff",
        2825 => x"631a350b",
        2826 => x"9307c000",
        2827 => x"2320f900",
        2828 => x"13050900",
        2829 => x"ef00401e",
        2830 => x"6f000001",
        2831 => x"e3d004fa",
        2832 => x"9307c000",
        2833 => x"2320f900",
        2834 => x"13050000",
        2835 => x"8320c101",
        2836 => x"03248101",
        2837 => x"83244101",
        2838 => x"03290101",
        2839 => x"8329c100",
        2840 => x"13010102",
        2841 => x"67800000",
        2842 => x"83270400",
        2843 => x"b3879740",
        2844 => x"63ce0704",
        2845 => x"1306b000",
        2846 => x"637af600",
        2847 => x"2320f400",
        2848 => x"3304f400",
        2849 => x"23209400",
        2850 => x"6f000001",
        2851 => x"83274400",
        2852 => x"631a8702",
        2853 => x"23a0f600",
        2854 => x"13050900",
        2855 => x"ef00c017",
        2856 => x"1305b400",
        2857 => x"93074400",
        2858 => x"137585ff",
        2859 => x"3307f540",
        2860 => x"e30ef5f8",
        2861 => x"3304e400",
        2862 => x"b387a740",
        2863 => x"2320f400",
        2864 => x"6ff0dff8",
        2865 => x"2322f700",
        2866 => x"6ff01ffd",
        2867 => x"13070400",
        2868 => x"03244400",
        2869 => x"6ff01ff2",
        2870 => x"13043500",
        2871 => x"1374c4ff",
        2872 => x"e30285fa",
        2873 => x"b305a440",
        2874 => x"13050900",
        2875 => x"ef00000e",
        2876 => x"e31a35f9",
        2877 => x"6ff05ff3",
        2878 => x"130101fe",
        2879 => x"232c8100",
        2880 => x"232e1100",
        2881 => x"232a9100",
        2882 => x"23282101",
        2883 => x"23263101",
        2884 => x"23244101",
        2885 => x"13040600",
        2886 => x"63940502",
        2887 => x"03248101",
        2888 => x"8320c101",
        2889 => x"83244101",
        2890 => x"03290101",
        2891 => x"8329c100",
        2892 => x"032a8100",
        2893 => x"93050600",
        2894 => x"13010102",
        2895 => x"6ff0dfe6",
        2896 => x"63180602",
        2897 => x"eff0dfd6",
        2898 => x"93040000",
        2899 => x"8320c101",
        2900 => x"03248101",
        2901 => x"03290101",
        2902 => x"8329c100",
        2903 => x"032a8100",
        2904 => x"13850400",
        2905 => x"83244101",
        2906 => x"13010102",
        2907 => x"67800000",
        2908 => x"130a0500",
        2909 => x"13890500",
        2910 => x"ef00400a",
        2911 => x"93090500",
        2912 => x"63688500",
        2913 => x"93571500",
        2914 => x"93040900",
        2915 => x"e3e087fc",
        2916 => x"93050400",
        2917 => x"13050a00",
        2918 => x"eff01fe1",
        2919 => x"93040500",
        2920 => x"e30605fa",
        2921 => x"13060400",
        2922 => x"63f48900",
        2923 => x"13860900",
        2924 => x"93050900",
        2925 => x"13850400",
        2926 => x"efe01fae",
        2927 => x"93050900",
        2928 => x"13050a00",
        2929 => x"eff0dfce",
        2930 => x"6ff05ff8",
        2931 => x"130101ff",
        2932 => x"23248100",
        2933 => x"23229100",
        2934 => x"13040500",
        2935 => x"13850500",
        2936 => x"23261100",
        2937 => x"23a20188",
        2938 => x"ef00000c",
        2939 => x"9307f0ff",
        2940 => x"6318f500",
        2941 => x"83a74188",
        2942 => x"63840700",
        2943 => x"2320f400",
        2944 => x"8320c100",
        2945 => x"03248100",
        2946 => x"83244100",
        2947 => x"13010101",
        2948 => x"67800000",
        2949 => x"67800000",
        2950 => x"67800000",
        2951 => x"83a7c5ff",
        2952 => x"1385c7ff",
        2953 => x"63d80700",
        2954 => x"b385a500",
        2955 => x"83a70500",
        2956 => x"3305f500",
        2957 => x"67800000",
        2958 => x"9308d005",
        2959 => x"73000000",
        2960 => x"63520502",
        2961 => x"130101ff",
        2962 => x"23248100",
        2963 => x"13040500",
        2964 => x"23261100",
        2965 => x"33048040",
        2966 => x"efe05fc6",
        2967 => x"23208500",
        2968 => x"6f000000",
        2969 => x"6f000000",
        2970 => x"130101ff",
        2971 => x"23261100",
        2972 => x"23248100",
        2973 => x"9308900a",
        2974 => x"73000000",
        2975 => x"13040500",
        2976 => x"635a0500",
        2977 => x"33048040",
        2978 => x"efe05fc3",
        2979 => x"23208500",
        2980 => x"1304f0ff",
        2981 => x"8320c100",
        2982 => x"13050400",
        2983 => x"03248100",
        2984 => x"13010101",
        2985 => x"67800000",
        2986 => x"83a70189",
        2987 => x"130101ff",
        2988 => x"23261100",
        2989 => x"93060500",
        2990 => x"13870189",
        2991 => x"639c0702",
        2992 => x"9308600d",
        2993 => x"13050000",
        2994 => x"73000000",
        2995 => x"9307f0ff",
        2996 => x"6310f502",
        2997 => x"efe09fbe",
        2998 => x"9307c000",
        2999 => x"2320f500",
        3000 => x"1305f0ff",
        3001 => x"8320c100",
        3002 => x"13010101",
        3003 => x"67800000",
        3004 => x"2320a700",
        3005 => x"83270700",
        3006 => x"9308600d",
        3007 => x"b386f600",
        3008 => x"13850600",
        3009 => x"73000000",
        3010 => x"e316d5fc",
        3011 => x"2320a700",
        3012 => x"13850700",
        3013 => x"6ff01ffd",
        3014 => x"10000000",
        3015 => x"00000000",
        3016 => x"037a5200",
        3017 => x"017c0101",
        3018 => x"1b0d0200",
        3019 => x"10000000",
        3020 => x"18000000",
        3021 => x"88d8ffff",
        3022 => x"78040000",
        3023 => x"00000000",
        3024 => x"10000000",
        3025 => x"00000000",
        3026 => x"037a5200",
        3027 => x"017c0101",
        3028 => x"1b0d0200",
        3029 => x"10000000",
        3030 => x"18000000",
        3031 => x"d8dcffff",
        3032 => x"50040000",
        3033 => x"00000000",
        3034 => x"10000000",
        3035 => x"00000000",
        3036 => x"037a5200",
        3037 => x"017c0101",
        3038 => x"1b0d0200",
        3039 => x"10000000",
        3040 => x"18000000",
        3041 => x"00e1ffff",
        3042 => x"30040000",
        3043 => x"00000000",
        3044 => x"10000000",
        3045 => x"00000000",
        3046 => x"037a5200",
        3047 => x"017c0101",
        3048 => x"1b0d0200",
        3049 => x"10000000",
        3050 => x"18000000",
        3051 => x"08e5ffff",
        3052 => x"e4030000",
        3053 => x"00000000",
        3054 => x"28020000",
        3055 => x"98010000",
        3056 => x"98010000",
        3057 => x"98010000",
        3058 => x"98010000",
        3059 => x"0c020000",
        3060 => x"98010000",
        3061 => x"cc010000",
        3062 => x"98010000",
        3063 => x"98010000",
        3064 => x"cc010000",
        3065 => x"98010000",
        3066 => x"98010000",
        3067 => x"98010000",
        3068 => x"98010000",
        3069 => x"98010000",
        3070 => x"98010000",
        3071 => x"98010000",
        3072 => x"7c010000",
        3073 => x"3c050000",
        3074 => x"24050000",
        3075 => x"24050000",
        3076 => x"24050000",
        3077 => x"24050000",
        3078 => x"54050000",
        3079 => x"a8050000",
        3080 => x"d0050000",
        3081 => x"24050000",
        3082 => x"24050000",
        3083 => x"24050000",
        3084 => x"24050000",
        3085 => x"24050000",
        3086 => x"24050000",
        3087 => x"24050000",
        3088 => x"24050000",
        3089 => x"24050000",
        3090 => x"24050000",
        3091 => x"24050000",
        3092 => x"24050000",
        3093 => x"24050000",
        3094 => x"24050000",
        3095 => x"c4040000",
        3096 => x"c4040000",
        3097 => x"24050000",
        3098 => x"24050000",
        3099 => x"24050000",
        3100 => x"24050000",
        3101 => x"24050000",
        3102 => x"24050000",
        3103 => x"24050000",
        3104 => x"24050000",
        3105 => x"24050000",
        3106 => x"24050000",
        3107 => x"24050000",
        3108 => x"24050000",
        3109 => x"54050000",
        3110 => x"3c050000",
        3111 => x"78050000",
        3112 => x"90050000",
        3113 => x"24050000",
        3114 => x"24050000",
        3115 => x"24050000",
        3116 => x"24050000",
        3117 => x"24050000",
        3118 => x"24050000",
        3119 => x"60050000",
        3120 => x"24050000",
        3121 => x"24050000",
        3122 => x"24050000",
        3123 => x"24050000",
        3124 => x"c4040000",
        3125 => x"c4040000",
        3126 => x"00010202",
        3127 => x"03030303",
        3128 => x"04040404",
        3129 => x"04040404",
        3130 => x"05050505",
        3131 => x"05050505",
        3132 => x"05050505",
        3133 => x"05050505",
        3134 => x"06060606",
        3135 => x"06060606",
        3136 => x"06060606",
        3137 => x"06060606",
        3138 => x"06060606",
        3139 => x"06060606",
        3140 => x"06060606",
        3141 => x"06060606",
        3142 => x"07070707",
        3143 => x"07070707",
        3144 => x"07070707",
        3145 => x"07070707",
        3146 => x"07070707",
        3147 => x"07070707",
        3148 => x"07070707",
        3149 => x"07070707",
        3150 => x"07070707",
        3151 => x"07070707",
        3152 => x"07070707",
        3153 => x"07070707",
        3154 => x"07070707",
        3155 => x"07070707",
        3156 => x"07070707",
        3157 => x"07070707",
        3158 => x"08080808",
        3159 => x"08080808",
        3160 => x"08080808",
        3161 => x"08080808",
        3162 => x"08080808",
        3163 => x"08080808",
        3164 => x"08080808",
        3165 => x"08080808",
        3166 => x"08080808",
        3167 => x"08080808",
        3168 => x"08080808",
        3169 => x"08080808",
        3170 => x"08080808",
        3171 => x"08080808",
        3172 => x"08080808",
        3173 => x"08080808",
        3174 => x"08080808",
        3175 => x"08080808",
        3176 => x"08080808",
        3177 => x"08080808",
        3178 => x"08080808",
        3179 => x"08080808",
        3180 => x"08080808",
        3181 => x"08080808",
        3182 => x"08080808",
        3183 => x"08080808",
        3184 => x"08080808",
        3185 => x"08080808",
        3186 => x"08080808",
        3187 => x"08080808",
        3188 => x"08080808",
        3189 => x"08080808",
        3190 => x"0d0a0d0a",
        3191 => x"44697370",
        3192 => x"6c617969",
        3193 => x"6e672074",
        3194 => x"68652074",
        3195 => x"696d6520",
        3196 => x"70617373",
        3197 => x"65642073",
        3198 => x"696e6365",
        3199 => x"20726573",
        3200 => x"65740d0a",
        3201 => x"0d0a0000",
        3202 => x"2530356c",
        3203 => x"643a2530",
        3204 => x"366c6420",
        3205 => x"20202530",
        3206 => x"326c643a",
        3207 => x"2530326c",
        3208 => x"643a2530",
        3209 => x"326c640d",
        3210 => x"00000000",
        3211 => x"696e7465",
        3212 => x"72727570",
        3213 => x"74000000",
        3214 => x"52495343",
        3215 => x"2d562052",
        3216 => x"56333249",
        3217 => x"4d206261",
        3218 => x"7265206d",
        3219 => x"6574616c",
        3220 => x"2070726f",
        3221 => x"63657373",
        3222 => x"6f720000",
        3223 => x"54686520",
        3224 => x"48616775",
        3225 => x"6520556e",
        3226 => x"69766572",
        3227 => x"73697479",
        3228 => x"206f6620",
        3229 => x"4170706c",
        3230 => x"69656420",
        3231 => x"53636965",
        3232 => x"6e636573",
        3233 => x"00000000",
        3234 => x"44657061",
        3235 => x"72746d65",
        3236 => x"6e74206f",
        3237 => x"6620456c",
        3238 => x"65637472",
        3239 => x"6963616c",
        3240 => x"20456e67",
        3241 => x"696e6565",
        3242 => x"72696e67",
        3243 => x"00000000",
        3244 => x"4a2e452e",
        3245 => x"4a2e206f",
        3246 => x"70206465",
        3247 => x"6e204272",
        3248 => x"6f757700",
        3249 => x"3c627265",
        3250 => x"616b3e0d",
        3251 => x"0a000000",
        3252 => x"0d0a4542",
        3253 => x"5245414b",
        3254 => x"21206d69",
        3255 => x"70203d20",
        3256 => x"00000000",
        3257 => x"232d302b",
        3258 => x"20000000",
        3259 => x"686c4c00",
        3260 => x"65666745",
        3261 => x"46470000",
        3262 => x"30313233",
        3263 => x"34353637",
        3264 => x"38394142",
        3265 => x"43444546",
        3266 => x"00000000",
        3267 => x"30313233",
        3268 => x"34353637",
        3269 => x"38396162",
        3270 => x"63646566",
        3271 => x"00000000",
        3272 => x"dc250000",
        3273 => x"fc250000",
        3274 => x"a8250000",
        3275 => x"a8250000",
        3276 => x"a8250000",
        3277 => x"a8250000",
        3278 => x"fc250000",
        3279 => x"a8250000",
        3280 => x"a8250000",
        3281 => x"a8250000",
        3282 => x"a8250000",
        3283 => x"e8270000",
        3284 => x"54260000",
        3285 => x"64270000",
        3286 => x"a8250000",
        3287 => x"a8250000",
        3288 => x"30280000",
        3289 => x"a8250000",
        3290 => x"54260000",
        3291 => x"a8250000",
        3292 => x"a8250000",
        3293 => x"70270000",
        3294 => x"18000020",
        3295 => x"2c320000",
        3296 => x"38320000",
        3297 => x"5c320000",
        3298 => x"88320000",
        3299 => x"b0320000",
        3300 => x"00000000",
        3301 => x"00000000",
        3302 => x"00000000",
        3303 => x"00000000",
        3304 => x"00000000",
        3305 => x"00000000",
        3306 => x"00000000",
        3307 => x"00000000",
        3308 => x"00000000",
        3309 => x"00000000",
        3310 => x"00000000",
        3311 => x"00000000",
        3312 => x"00000000",
        3313 => x"00000000",
        3314 => x"00000000",
        3315 => x"00000000",
        3316 => x"00000000",
        3317 => x"00000000",
        3318 => x"00000000",
        3319 => x"00000000",
        3320 => x"00000000",
        3321 => x"00000000",
        3322 => x"00000000",
        3323 => x"00000000",
        3324 => x"00000000",
        3325 => x"80000020",
        3326 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
