-- srec2vhdl table generator
-- for input file flash.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97",    1 => x"11",    2 => x"00",    3 => x"20", 
           4 => x"93",    5 => x"81",    6 => x"01",    7 => x"81", 
           8 => x"17",    9 => x"41",   10 => x"00",   11 => x"20", 
          12 => x"13",   13 => x"01",   14 => x"81",   15 => x"ff", 
          16 => x"97",   17 => x"00",   18 => x"00",   19 => x"00", 
          20 => x"e7",   21 => x"80",   22 => x"c0",   23 => x"00", 
          24 => x"6f",   25 => x"00",   26 => x"00",   27 => x"00", 
          28 => x"13",   29 => x"01",   30 => x"01",   31 => x"fe", 
          32 => x"23",   33 => x"2e",   34 => x"81",   35 => x"00", 
          36 => x"13",   37 => x"04",   38 => x"01",   39 => x"02", 
          40 => x"b7",   41 => x"07",   42 => x"00",   43 => x"f0", 
          44 => x"93",   45 => x"87",   46 => x"47",   47 => x"00", 
          48 => x"23",   49 => x"26",   50 => x"f4",   51 => x"fe", 
          52 => x"b7",   53 => x"07",   54 => x"00",   55 => x"20", 
          56 => x"83",   57 => x"a7",   58 => x"07",   59 => x"00", 
          60 => x"13",   61 => x"87",   62 => x"17",   63 => x"00", 
          64 => x"b7",   65 => x"07",   66 => x"00",   67 => x"20", 
          68 => x"23",   69 => x"a0",   70 => x"e7",   71 => x"00", 
          72 => x"23",   73 => x"24",   74 => x"04",   75 => x"fe", 
          76 => x"6f",   77 => x"00",   78 => x"00",   79 => x"01", 
          80 => x"83",   81 => x"27",   82 => x"84",   83 => x"fe", 
          84 => x"93",   85 => x"87",   86 => x"17",   87 => x"00", 
          88 => x"23",   89 => x"24",   90 => x"f4",   91 => x"fe", 
          92 => x"03",   93 => x"27",   94 => x"84",   95 => x"fe", 
          96 => x"b7",   97 => x"57",   98 => x"4c",   99 => x"00", 
         100 => x"93",  101 => x"87",  102 => x"f7",  103 => x"b3", 
         104 => x"e3",  105 => x"f4",  106 => x"e7",  107 => x"fe", 
         108 => x"83",  109 => x"27",  110 => x"c4",  111 => x"fe", 
         112 => x"13",  113 => x"07",  114 => x"f0",  115 => x"ff", 
         116 => x"23",  117 => x"a0",  118 => x"e7",  119 => x"00", 
         120 => x"23",  121 => x"24",  122 => x"04",  123 => x"fe", 
         124 => x"6f",  125 => x"00",  126 => x"00",  127 => x"01", 
         128 => x"83",  129 => x"27",  130 => x"84",  131 => x"fe", 
         132 => x"93",  133 => x"87",  134 => x"17",  135 => x"00", 
         136 => x"23",  137 => x"24",  138 => x"f4",  139 => x"fe", 
         140 => x"03",  141 => x"27",  142 => x"84",  143 => x"fe", 
         144 => x"b7",  145 => x"57",  146 => x"4c",  147 => x"00", 
         148 => x"93",  149 => x"87",  150 => x"f7",  151 => x"b3", 
         152 => x"e3",  153 => x"f4",  154 => x"e7",  155 => x"fe", 
         156 => x"83",  157 => x"27",  158 => x"c4",  159 => x"fe", 
         160 => x"23",  161 => x"a0",  162 => x"07",  163 => x"00", 
         164 => x"6f",  165 => x"f0",  166 => x"5f",  167 => x"fa", 
        others => (others => '-')
    );
end package processor_common_rom;
