--
-- This file is part of the THUAS RISC-V Minimal Project
--
-- (c)2022, Jesse E.J. op den Brouw <J.E.J.opdenBrouw@hhs.nl>
--
-- bootloader.vhd - Description of the bootloader ROM unit

-- This hardware description is for educational purposes only. 
-- This hardware description is distributed in the hope that it
-- will be useful, but WITHOUT ANY WARRANTY; without even the
-- implied warranty of MERCHANTABILITY or FITNESS FOR A
-- PARTICULAR PURPOSE.

-- This file contains the description of the boot ROM. The ROM
-- is placed in immutable onboard RAM blocks. A read takes two
-- clock cycles, for both instruction and data.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.processor_common.all;
use work.processor_common_rom.all;

entity bootloader is
    port (I_clk : in std_logic;
          I_areset : in std_logic;
          I_pc : in data_type;
          I_address : in data_type;
          I_csboot : in std_logic;
          I_size : in size_type;
          I_stall : in std_logic;
          O_instr : out data_type;
          O_data_out : out data_type;
          --
          O_instruction_misaligned_error : out std_logic;
          O_load_misaligned_error : out std_logic
         );
end entity bootloader;

architecture rtl of bootloader is

-- The bootloader ROM
signal bootrom : bootloader_type := (
           0 => x"97110010",
           1 => x"93810180",
           2 => x"17810010",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"9382c23c",
           6 => x"73905230",
           7 => x"b7070020",
           8 => x"37050020",
           9 => x"93870700",
          10 => x"13070500",
          11 => x"13060000",
          12 => x"63e4e700",
          13 => x"3386e740",
          14 => x"93050000",
          15 => x"13050500",
          16 => x"ef00403c",
          17 => x"37050020",
          18 => x"b7070020",
          19 => x"93870700",
          20 => x"13070500",
          21 => x"13060000",
          22 => x"63e4e700",
          23 => x"3386e740",
          24 => x"b7150010",
          25 => x"938585bb",
          26 => x"13050500",
          27 => x"ef004037",
          28 => x"ef00003d",
          29 => x"6f000000",
          30 => x"37170000",
          31 => x"b70700f0",
          32 => x"13077745",
          33 => x"23a2e702",
          34 => x"67800000",
          35 => x"1375f50f",
          36 => x"b70700f0",
          37 => x"23a0a702",
          38 => x"370700f0",
          39 => x"8327c702",
          40 => x"93f70701",
          41 => x"e38c07fe",
          42 => x"67800000",
          43 => x"130101ff",
          44 => x"23248100",
          45 => x"23261100",
          46 => x"13040500",
          47 => x"03450400",
          48 => x"631a0500",
          49 => x"8320c100",
          50 => x"03248100",
          51 => x"13010101",
          52 => x"67800000",
          53 => x"13041400",
          54 => x"eff05ffb",
          55 => x"6ff01ffe",
          56 => x"63040500",
          57 => x"6ff09ffc",
          58 => x"67800000",
          59 => x"b70600f0",
          60 => x"83a7c602",
          61 => x"93f74700",
          62 => x"e38c07fe",
          63 => x"03a50602",
          64 => x"1375f50f",
          65 => x"67800000",
          66 => x"b70700f0",
          67 => x"03a5c702",
          68 => x"13754500",
          69 => x"67800000",
          70 => x"130101fd",
          71 => x"23248102",
          72 => x"23229102",
          73 => x"23202103",
          74 => x"232e3101",
          75 => x"232c4101",
          76 => x"232a5101",
          77 => x"23286101",
          78 => x"23267101",
          79 => x"23248101",
          80 => x"23229101",
          81 => x"23261102",
          82 => x"93040500",
          83 => x"13040000",
          84 => x"9309d000",
          85 => x"1389f5ff",
          86 => x"130ae005",
          87 => x"930a5001",
          88 => x"130b8000",
          89 => x"930ba000",
          90 => x"130c3000",
          91 => x"b71c0010",
          92 => x"eff0dff7",
          93 => x"93070500",
          94 => x"1375f50f",
          95 => x"63043509",
          96 => x"63cca902",
          97 => x"63006505",
          98 => x"630e7507",
          99 => x"63008507",
         100 => x"63562407",
         101 => x"93f7f70f",
         102 => x"138707fe",
         103 => x"1377f70f",
         104 => x"e368eafc",
         105 => x"33878400",
         106 => x"2300f700",
         107 => x"13041400",
         108 => x"eff0dfed",
         109 => x"6ff0dffb",
         110 => x"63065503",
         111 => x"1307f007",
         112 => x"e318e5fc",
         113 => x"630c0402",
         114 => x"1305f007",
         115 => x"eff01fec",
         116 => x"1304f4ff",
         117 => x"6ff0dff9",
         118 => x"1305f007",
         119 => x"eff01feb",
         120 => x"1304f4ff",
         121 => x"e31a04fe",
         122 => x"6ff09ff8",
         123 => x"13858caa",
         124 => x"eff0dfeb",
         125 => x"13040000",
         126 => x"6ff09ff7",
         127 => x"13057000",
         128 => x"6ff01ffb",
         129 => x"b3848400",
         130 => x"37150010",
         131 => x"23800400",
         132 => x"13050598",
         133 => x"eff09fe9",
         134 => x"8320c102",
         135 => x"13050400",
         136 => x"03248102",
         137 => x"83244102",
         138 => x"03290102",
         139 => x"8329c101",
         140 => x"032a8101",
         141 => x"832a4101",
         142 => x"032b0101",
         143 => x"832bc100",
         144 => x"032c8100",
         145 => x"832c4100",
         146 => x"13010103",
         147 => x"67800000",
         148 => x"37180010",
         149 => x"93070500",
         150 => x"130858ab",
         151 => x"03c70700",
         152 => x"33070701",
         153 => x"03470700",
         154 => x"13778700",
         155 => x"63160702",
         156 => x"13050000",
         157 => x"93081000",
         158 => x"83c60700",
         159 => x"3307d800",
         160 => x"03470700",
         161 => x"13764704",
         162 => x"631c0600",
         163 => x"63840500",
         164 => x"23a0f500",
         165 => x"67800000",
         166 => x"93871700",
         167 => x"6ff01ffc",
         168 => x"13734700",
         169 => x"13154500",
         170 => x"13860600",
         171 => x"630a0300",
         172 => x"938606fd",
         173 => x"33e5a600",
         174 => x"93871700",
         175 => x"6ff0dffb",
         176 => x"13773700",
         177 => x"63141701",
         178 => x"13860602",
         179 => x"130696fa",
         180 => x"3365a600",
         181 => x"6ff05ffe",
         182 => x"130101fe",
         183 => x"232e1100",
         184 => x"23220100",
         185 => x"23240100",
         186 => x"23060100",
         187 => x"9386f5ff",
         188 => x"13077000",
         189 => x"93070500",
         190 => x"6374d700",
         191 => x"93058000",
         192 => x"13054100",
         193 => x"b305b500",
         194 => x"13069003",
         195 => x"93f6f700",
         196 => x"13870603",
         197 => x"6374e600",
         198 => x"13877605",
         199 => x"a38fe5fe",
         200 => x"9385f5ff",
         201 => x"93d74700",
         202 => x"e312b5fe",
         203 => x"eff05fdb",
         204 => x"8320c101",
         205 => x"13010102",
         206 => x"67800000",
         207 => x"130101fe",
         208 => x"23263101",
         209 => x"b7190010",
         210 => x"232c8100",
         211 => x"232a9100",
         212 => x"23282101",
         213 => x"23244101",
         214 => x"232e1100",
         215 => x"93040500",
         216 => x"13090000",
         217 => x"13040000",
         218 => x"938959ab",
         219 => x"130a1000",
         220 => x"63449902",
         221 => x"8320c101",
         222 => x"13050400",
         223 => x"03248101",
         224 => x"83244101",
         225 => x"03290101",
         226 => x"8329c100",
         227 => x"032a8100",
         228 => x"13010102",
         229 => x"67800000",
         230 => x"eff05fd5",
         231 => x"b3073501",
         232 => x"83c70700",
         233 => x"13144400",
         234 => x"13f74700",
         235 => x"630a0700",
         236 => x"930705fd",
         237 => x"3364f400",
         238 => x"13091900",
         239 => x"6ff05ffb",
         240 => x"13f74704",
         241 => x"e30a07fe",
         242 => x"93f73700",
         243 => x"63944701",
         244 => x"13050502",
         245 => x"930795fa",
         246 => x"6ff0dffd",
         247 => x"6f000000",
         248 => x"13030500",
         249 => x"630e0600",
         250 => x"83830500",
         251 => x"23007300",
         252 => x"1306f6ff",
         253 => x"13031300",
         254 => x"93851500",
         255 => x"e31606fe",
         256 => x"67800000",
         257 => x"13030500",
         258 => x"630a0600",
         259 => x"2300b300",
         260 => x"1306f6ff",
         261 => x"13031300",
         262 => x"e31a06fe",
         263 => x"67800000",
         264 => x"03460500",
         265 => x"83c60500",
         266 => x"13051500",
         267 => x"93851500",
         268 => x"6314d600",
         269 => x"e31606fe",
         270 => x"3305d640",
         271 => x"67800000",
         272 => x"130101f8",
         273 => x"232e1106",
         274 => x"232c8106",
         275 => x"232a9106",
         276 => x"23282107",
         277 => x"23263107",
         278 => x"23244107",
         279 => x"23225107",
         280 => x"23206107",
         281 => x"232e7105",
         282 => x"232c8105",
         283 => x"232a9105",
         284 => x"2328a105",
         285 => x"2326b105",
         286 => x"eff01fc0",
         287 => x"37150010",
         288 => x"13058595",
         289 => x"eff0dfc5",
         290 => x"b70700f0",
         291 => x"1307f03f",
         292 => x"b704a000",
         293 => x"37091000",
         294 => x"23a2e700",
         295 => x"13041000",
         296 => x"93841400",
         297 => x"1309f9ff",
         298 => x"b70900f0",
         299 => x"eff0dfc5",
         300 => x"631a050e",
         301 => x"13041400",
         302 => x"6316940c",
         303 => x"b70700f0",
         304 => x"23a20700",
         305 => x"63140500",
         306 => x"e7000500",
         307 => x"eff01fc2",
         308 => x"93071002",
         309 => x"93040000",
         310 => x"6316f520",
         311 => x"371b0010",
         312 => x"1305cb97",
         313 => x"b70901ff",
         314 => x"370a0001",
         315 => x"b70affff",
         316 => x"eff01fbf",
         317 => x"9389f9ff",
         318 => x"130afaff",
         319 => x"938afa0f",
         320 => x"370400f0",
         321 => x"83274400",
         322 => x"93c71700",
         323 => x"2322f400",
         324 => x"eff0dfbd",
         325 => x"1375f50f",
         326 => x"93073005",
         327 => x"6314f51a",
         328 => x"eff0dfbc",
         329 => x"1374f50f",
         330 => x"9307f4fc",
         331 => x"93f7f70f",
         332 => x"13072000",
         333 => x"6368f712",
         334 => x"93071003",
         335 => x"6318f406",
         336 => x"13052000",
         337 => x"eff09fdf",
         338 => x"1309d5ff",
         339 => x"13054000",
         340 => x"eff0dfde",
         341 => x"13040500",
         342 => x"3309a900",
         343 => x"130c3000",
         344 => x"930c1000",
         345 => x"631a2407",
         346 => x"1304a000",
         347 => x"eff01fb8",
         348 => x"1375f50f",
         349 => x"e31c85fe",
         350 => x"1305cb97",
         351 => x"eff05fb6",
         352 => x"6ff01ff8",
         353 => x"b3772401",
         354 => x"e39207f2",
         355 => x"1305a002",
         356 => x"eff0dfaf",
         357 => x"83a74900",
         358 => x"93d71700",
         359 => x"23a2f900",
         360 => x"6ff0dff0",
         361 => x"13051000",
         362 => x"6ff05ff1",
         363 => x"93072003",
         364 => x"13052000",
         365 => x"631af400",
         366 => x"eff05fd8",
         367 => x"1309c5ff",
         368 => x"13056000",
         369 => x"6ff0dff8",
         370 => x"eff05fd7",
         371 => x"1309b5ff",
         372 => x"13058000",
         373 => x"6ff0dff7",
         374 => x"13052000",
         375 => x"eff01fd6",
         376 => x"2324a100",
         377 => x"937bc4ff",
         378 => x"83a70b00",
         379 => x"13072000",
         380 => x"2326f100",
         381 => x"93773400",
         382 => x"6382e704",
         383 => x"638a8705",
         384 => x"63849703",
         385 => x"8327c100",
         386 => x"03278100",
         387 => x"93f707f0",
         388 => x"b3e7e700",
         389 => x"2326f100",
         390 => x"8327c100",
         391 => x"13041400",
         392 => x"23a0fb00",
         393 => x"6ff01ff4",
         394 => x"8327c100",
         395 => x"03278100",
         396 => x"b3f75701",
         397 => x"13178700",
         398 => x"6ff09ffd",
         399 => x"8327c100",
         400 => x"03278100",
         401 => x"b3f73701",
         402 => x"13170701",
         403 => x"6ff05ffc",
         404 => x"8327c100",
         405 => x"03278100",
         406 => x"b3f74701",
         407 => x"13178701",
         408 => x"6ff01ffb",
         409 => x"930794fc",
         410 => x"93f7f70f",
         411 => x"1309a000",
         412 => x"6362f704",
         413 => x"13052000",
         414 => x"eff05fcc",
         415 => x"93077003",
         416 => x"13058000",
         417 => x"630af400",
         418 => x"93078003",
         419 => x"13056000",
         420 => x"6304f400",
         421 => x"13054000",
         422 => x"eff05fca",
         423 => x"93040500",
         424 => x"1304a000",
         425 => x"eff09fa4",
         426 => x"1375f50f",
         427 => x"e31c85fe",
         428 => x"6ff09fec",
         429 => x"eff09fa3",
         430 => x"1375f50f",
         431 => x"e31c25ff",
         432 => x"6ff09feb",
         433 => x"9307a004",
         434 => x"6310f508",
         435 => x"23220402",
         436 => x"23220400",
         437 => x"e7800400",
         438 => x"b70700f0",
         439 => x"1307a00a",
         440 => x"23a2e700",
         441 => x"37190010",
         442 => x"13050998",
         443 => x"b7190010",
         444 => x"eff01f9f",
         445 => x"13040000",
         446 => x"b71b0010",
         447 => x"938959ab",
         448 => x"b7170010",
         449 => x"13854798",
         450 => x"eff09f9d",
         451 => x"93059002",
         452 => x"13054101",
         453 => x"eff05fa0",
         454 => x"13054101",
         455 => x"ef00401e",
         456 => x"b7170010",
         457 => x"130a0500",
         458 => x"93858798",
         459 => x"13054101",
         460 => x"eff01fcf",
         461 => x"63100502",
         462 => x"37150010",
         463 => x"1305c598",
         464 => x"eff01f9a",
         465 => x"6f004003",
         466 => x"93073002",
         467 => x"e316f5e2",
         468 => x"6ff09ff8",
         469 => x"b7170010",
         470 => x"938547a7",
         471 => x"13054101",
         472 => x"eff01fcc",
         473 => x"63100502",
         474 => x"b70700f0",
         475 => x"23a20702",
         476 => x"23a20700",
         477 => x"e7800400",
         478 => x"13050998",
         479 => x"eff05f96",
         480 => x"6ff01ff8",
         481 => x"b7170010",
         482 => x"13063000",
         483 => x"938587a7",
         484 => x"13054101",
         485 => x"ef008018",
         486 => x"63100504",
         487 => x"93050000",
         488 => x"13057101",
         489 => x"eff0dfaa",
         490 => x"93773500",
         491 => x"13040500",
         492 => x"639a0712",
         493 => x"93058000",
         494 => x"eff01fb2",
         495 => x"37150010",
         496 => x"1305c5a7",
         497 => x"eff0df91",
         498 => x"03250400",
         499 => x"93058000",
         500 => x"eff09fb0",
         501 => x"6ff05ffa",
         502 => x"b7170010",
         503 => x"13063000",
         504 => x"938587a9",
         505 => x"13054101",
         506 => x"ef004013",
         507 => x"63180502",
         508 => x"93050101",
         509 => x"13057101",
         510 => x"eff09fa5",
         511 => x"93773500",
         512 => x"13040500",
         513 => x"6390070e",
         514 => x"03250101",
         515 => x"93050000",
         516 => x"eff01fa4",
         517 => x"2320a400",
         518 => x"6ff01ff6",
         519 => x"13063000",
         520 => x"9385cba9",
         521 => x"13054101",
         522 => x"ef00400f",
         523 => x"83474101",
         524 => x"1307e006",
         525 => x"63080508",
         526 => x"639ce70a",
         527 => x"93773400",
         528 => x"6392070a",
         529 => x"130c0404",
         530 => x"b71c0010",
         531 => x"371d0010",
         532 => x"930d80ff",
         533 => x"93058000",
         534 => x"13050400",
         535 => x"eff0dfa7",
         536 => x"1385cca7",
         537 => x"eff0df87",
         538 => x"032a0400",
         539 => x"93058000",
         540 => x"930a8001",
         541 => x"13050a00",
         542 => x"eff01fa6",
         543 => x"13050daa",
         544 => x"eff01f86",
         545 => x"370b00ff",
         546 => x"33756a01",
         547 => x"33555501",
         548 => x"b3063501",
         549 => x"83c60600",
         550 => x"93f67609",
         551 => x"63800604",
         552 => x"938a8aff",
         553 => x"eff08ffe",
         554 => x"135b8b00",
         555 => x"e39ebafd",
         556 => x"13044400",
         557 => x"13050998",
         558 => x"eff09f82",
         559 => x"e31c8cf8",
         560 => x"6ff09feb",
         561 => x"e38ce7f6",
         562 => x"93050000",
         563 => x"13057101",
         564 => x"eff01f98",
         565 => x"13040500",
         566 => x"6ff05ff6",
         567 => x"1305e002",
         568 => x"6ff01ffc",
         569 => x"37150010",
         570 => x"130505a8",
         571 => x"6ff05fe5",
         572 => x"e3040ae8",
         573 => x"37150010",
         574 => x"130545aa",
         575 => x"6ff05fe4",
         576 => x"93070500",
         577 => x"03c70700",
         578 => x"93871700",
         579 => x"e31c07fe",
         580 => x"3385a740",
         581 => x"1305f5ff",
         582 => x"67800000",
         583 => x"630a0602",
         584 => x"1306f6ff",
         585 => x"13070000",
         586 => x"b307e500",
         587 => x"b386e500",
         588 => x"83c70700",
         589 => x"83c60600",
         590 => x"6398d700",
         591 => x"6306c700",
         592 => x"13071700",
         593 => x"e39207fe",
         594 => x"3385d740",
         595 => x"67800000",
         596 => x"13050000",
         597 => x"67800000",
         598 => x"0d0a5448",
         599 => x"55415320",
         600 => x"52495343",
         601 => x"2d562042",
         602 => x"6f6f746c",
         603 => x"6f616465",
         604 => x"72207630",
         605 => x"2e310d0a",
         606 => x"00000000",
         607 => x"3f0a0000",
         608 => x"0d0a0000",
         609 => x"3e200000",
         610 => x"68000000",
         611 => x"48656c70",
         612 => x"3a0d0a20",
         613 => x"68202020",
         614 => x"20202020",
         615 => x"20202020",
         616 => x"20202020",
         617 => x"202d2074",
         618 => x"68697320",
         619 => x"68656c70",
         620 => x"0d0a2072",
         621 => x"20202020",
         622 => x"20202020",
         623 => x"20202020",
         624 => x"20202020",
         625 => x"2d207275",
         626 => x"6e206170",
         627 => x"706c6963",
         628 => x"6174696f",
         629 => x"6e0d0a20",
         630 => x"7277203c",
         631 => x"61646472",
         632 => x"3e202020",
         633 => x"20202020",
         634 => x"202d2072",
         635 => x"65616420",
         636 => x"776f7264",
         637 => x"2066726f",
         638 => x"6d206164",
         639 => x"64720d0a",
         640 => x"20777720",
         641 => x"3c616464",
         642 => x"723e203c",
         643 => x"64617461",
         644 => x"3e202d20",
         645 => x"77726974",
         646 => x"65206461",
         647 => x"74612061",
         648 => x"74206164",
         649 => x"64720d0a",
         650 => x"20647720",
         651 => x"3c616464",
         652 => x"723e2020",
         653 => x"20202020",
         654 => x"20202d20",
         655 => x"64756d70",
         656 => x"20313620",
         657 => x"776f7264",
         658 => x"730d0a20",
         659 => x"6e202020",
         660 => x"20202020",
         661 => x"20202020",
         662 => x"20202020",
         663 => x"202d2064",
         664 => x"756d7020",
         665 => x"6e657874",
         666 => x"20313620",
         667 => x"776f7264",
         668 => x"73000000",
         669 => x"72000000",
         670 => x"72772000",
         671 => x"3a200000",
         672 => x"4e6f7420",
         673 => x"6f6e2034",
         674 => x"2d627974",
         675 => x"6520626f",
         676 => x"756e6461",
         677 => x"72792100",
         678 => x"77772000",
         679 => x"64772000",
         680 => x"20200000",
         681 => x"3f3f0000",
         682 => x"3c627265",
         683 => x"616b3e0d",
         684 => x"0a000000",
         685 => x"00202020",
         686 => x"20202020",
         687 => x"20202828",
         688 => x"28282820",
         689 => x"20202020",
         690 => x"20202020",
         691 => x"20202020",
         692 => x"20202020",
         693 => x"20881010",
         694 => x"10101010",
         695 => x"10101010",
         696 => x"10101010",
         697 => x"10040404",
         698 => x"04040404",
         699 => x"04040410",
         700 => x"10101010",
         701 => x"10104141",
         702 => x"41414141",
         703 => x"01010101",
         704 => x"01010101",
         705 => x"01010101",
         706 => x"01010101",
         707 => x"01010101",
         708 => x"10101010",
         709 => x"10104242",
         710 => x"42424242",
         711 => x"02020202",
         712 => x"02020202",
         713 => x"02020202",
         714 => x"02020202",
         715 => x"02020202",
         716 => x"10101010",
         717 => x"20000000",
         718 => x"00000000",
         719 => x"00000000",
         720 => x"00000000",
         721 => x"00000000",
         722 => x"00000000",
         723 => x"00000000",
         724 => x"00000000",
         725 => x"00000000",
         726 => x"00000000",
         727 => x"00000000",
         728 => x"00000000",
         729 => x"00000000",
         730 => x"00000000",
         731 => x"00000000",
         732 => x"00000000",
         733 => x"00000000",
         734 => x"00000000",
         735 => x"00000000",
         736 => x"00000000",
         737 => x"00000000",
         738 => x"00000000",
         739 => x"00000000",
         740 => x"00000000",
         741 => x"00000000",
         742 => x"00000000",
         743 => x"00000000",
         744 => x"00000000",
         745 => x"00000000",
         746 => x"00000000",
         747 => x"00000000",
         748 => x"00000000",
         749 => x"00000000",
         others => (others => '0')
        );

begin

    gen_bootrom: if HAVE_BOOT_ROM generate
        O_instruction_misaligned_error <= '0' when I_pc(1 downto 0) = "00" else '1';        

        -- ROM, for both instructions and read-only data
        process (I_clk, I_areset, I_pc, I_address, I_csboot, I_size, I_stall) is
        variable address_instr : integer range 0 to bootloader_size-1;
        variable address_data : integer range 0 to bootloader_size-1;
        variable instr_var : data_type;
        variable instr_recode : data_type;
        variable romdata_var : data_type;
        constant x : data_type := (others => 'X');
        begin
            -- Calculate addresses
            address_instr := to_integer(unsigned(I_pc(bootloader_size_bits-1 downto 2)));
            address_data := to_integer(unsigned(I_address(bootloader_size_bits-1 downto 2)));

            -- Quartus will detect ROM table and uses onboard RAM
            -- Do not use reset, otherwise ROM will be created with ALMs
            if rising_edge(I_clk) then
                if I_stall = '0' then
                    instr_var := bootrom(address_instr);
                end if;
                romdata_var := bootrom(address_data);
            end if;
            
            -- Recode instruction
            O_instr <= instr_var(7 downto 0) & instr_var(15 downto 8) & instr_var(23 downto 16) & instr_var(31 downto 24);
            
            O_load_misaligned_error <= '0';
            
            -- By natural size, for data
            if I_csboot = '1' then
                if I_size = size_word and I_address(1 downto 0) = "00" then
                    O_data_out <= romdata_var(7 downto 0) & romdata_var(15 downto 8) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_size = size_halfword and I_address(1 downto 0) = "00" then
                    O_data_out <= x(31 downto 16) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_size = size_halfword and I_address(1 downto 0) = "10" then
                    O_data_out <= x(31 downto 16) & romdata_var(7 downto 0) & romdata_var(15 downto 8);
                elsif I_size = size_byte then
                    case I_address(1 downto 0) is
                        when "00" => O_data_out <= x(31 downto 8) & romdata_var(31 downto 24);
                        when "01" => O_data_out <= x(31 downto 8) & romdata_var(23 downto 16);
                        when "10" => O_data_out <= x(31 downto 8) & romdata_var(15 downto 8);
                        when "11" => O_data_out <= x(31 downto 8) & romdata_var(7 downto 0);
                        when others => O_data_out <= x; O_load_misaligned_error <= '1';
                    end case;
                else
                    -- Chip select, but not aligned
                    O_data_out <= x;
                    O_load_misaligned_error <= '1';
                end if;
            else
                -- No chip select, so no data
                O_data_out <= x;
            end if;
        end process;
    end generate;

    gen_bootrom_not: if not HAVE_BOOT_ROM generate
        O_instruction_misaligned_error <= '0';
        O_load_misaligned_error <= '0';
        O_data_out <= (others => 'X');
        O_instr  <= (others => 'X');
    end generate;
end architecture rtl;
