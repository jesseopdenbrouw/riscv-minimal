-- srec2vhdl table generator
-- for input file string.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"93",    1 => x"81",    2 => x"01",    3 => x"00", 
           4 => x"17",    5 => x"41",    6 => x"00",    7 => x"20", 
           8 => x"13",    9 => x"01",   10 => x"c1",   11 => x"ff", 
          12 => x"b7",   13 => x"07",   14 => x"00",   15 => x"20", 
          16 => x"93",   17 => x"80",   18 => x"47",   19 => x"06", 
          20 => x"b7",   21 => x"07",   22 => x"00",   23 => x"20", 
          24 => x"93",   25 => x"84",   26 => x"47",   27 => x"06", 
          28 => x"13",   29 => x"09",   30 => x"c0",   31 => x"28", 
          32 => x"6f",   33 => x"00",   34 => x"40",   35 => x"01", 
          36 => x"23",   37 => x"a0",   38 => x"00",   39 => x"00", 
          40 => x"93",   41 => x"87",   42 => x"00",   43 => x"00", 
          44 => x"93",   45 => x"80",   46 => x"47",   47 => x"00", 
          48 => x"83",   49 => x"a7",   50 => x"07",   51 => x"00", 
          52 => x"e3",   53 => x"e8",   54 => x"90",   55 => x"fe", 
          56 => x"b7",   57 => x"07",   58 => x"00",   59 => x"20", 
          60 => x"93",   61 => x"80",   62 => x"07",   63 => x"00", 
          64 => x"b7",   65 => x"07",   66 => x"00",   67 => x"20", 
          68 => x"93",   69 => x"84",   70 => x"07",   71 => x"06", 
          72 => x"6f",   73 => x"00",   74 => x"40",   75 => x"01", 
          76 => x"83",   77 => x"27",   78 => x"09",   79 => x"00", 
          80 => x"23",   81 => x"a0",   82 => x"f0",   83 => x"00", 
          84 => x"93",   85 => x"80",   86 => x"40",   87 => x"00", 
          88 => x"13",   89 => x"09",   90 => x"49",   91 => x"00", 
          92 => x"e3",   93 => x"e8",   94 => x"90",   95 => x"fe", 
          96 => x"ef",   97 => x"00",   98 => x"80",   99 => x"10", 
         100 => x"ef",  101 => x"00",  102 => x"c0",  103 => x"00", 
         104 => x"13",  105 => x"05",  106 => x"00",  107 => x"00", 
         108 => x"ef",  109 => x"00",  110 => x"00",  111 => x"0c", 
         112 => x"13",  113 => x"01",  114 => x"01",  115 => x"f7", 
         116 => x"23",  117 => x"26",  118 => x"11",  119 => x"08", 
         120 => x"23",  121 => x"24",  122 => x"81",  123 => x"08", 
         124 => x"13",  125 => x"04",  126 => x"01",  127 => x"09", 
         128 => x"93",  129 => x"07",  130 => x"00",  131 => x"27", 
         132 => x"03",  133 => x"a5",  134 => x"07",  135 => x"00", 
         136 => x"83",  137 => x"a5",  138 => x"47",  139 => x"00", 
         140 => x"03",  141 => x"a6",  142 => x"87",  143 => x"00", 
         144 => x"83",  145 => x"a6",  146 => x"c7",  147 => x"00", 
         148 => x"03",  149 => x"a7",  150 => x"07",  151 => x"01", 
         152 => x"83",  153 => x"a7",  154 => x"47",  155 => x"01", 
         156 => x"23",  157 => x"2c",  158 => x"a4",  159 => x"fc", 
         160 => x"23",  161 => x"2e",  162 => x"b4",  163 => x"fc", 
         164 => x"23",  165 => x"20",  166 => x"c4",  167 => x"fe", 
         168 => x"23",  169 => x"22",  170 => x"d4",  171 => x"fe", 
         172 => x"23",  173 => x"24",  174 => x"e4",  175 => x"fe", 
         176 => x"23",  177 => x"26",  178 => x"f4",  179 => x"fe", 
         180 => x"93",  181 => x"07",  182 => x"84",  183 => x"fd", 
         184 => x"13",  185 => x"85",  186 => x"07",  187 => x"00", 
         188 => x"ef",  189 => x"00",  190 => x"40",  191 => x"15", 
         192 => x"93",  193 => x"07",  194 => x"05",  195 => x"00", 
         196 => x"23",  197 => x"28",  198 => x"f4",  199 => x"f6", 
         200 => x"13",  201 => x"07",  202 => x"84",  203 => x"fd", 
         204 => x"93",  205 => x"07",  206 => x"44",  207 => x"f7", 
         208 => x"93",  209 => x"05",  210 => x"07",  211 => x"00", 
         212 => x"13",  213 => x"85",  214 => x"07",  215 => x"00", 
         216 => x"ef",  217 => x"00",  218 => x"c0",  219 => x"11", 
         220 => x"93",  221 => x"07",  222 => x"84",  223 => x"fd", 
         224 => x"93",  225 => x"85",  226 => x"07",  227 => x"00", 
         228 => x"13",  229 => x"05",  230 => x"80",  231 => x"26", 
         232 => x"ef",  233 => x"00",  234 => x"40",  235 => x"02", 
         236 => x"93",  237 => x"07",  238 => x"05",  239 => x"00", 
         240 => x"23",  241 => x"28",  242 => x"f4",  243 => x"f6", 
         244 => x"83",  245 => x"27",  246 => x"04",  247 => x"f7", 
         248 => x"13",  249 => x"85",  250 => x"07",  251 => x"00", 
         252 => x"83",  253 => x"20",  254 => x"c1",  255 => x"08", 
         256 => x"03",  257 => x"24",  258 => x"81",  259 => x"08", 
         260 => x"13",  261 => x"01",  262 => x"01",  263 => x"09", 
         264 => x"67",  265 => x"80",  266 => x"00",  267 => x"00", 
         268 => x"03",  269 => x"46",  270 => x"05",  271 => x"00", 
         272 => x"83",  273 => x"c6",  274 => x"05",  275 => x"00", 
         276 => x"13",  277 => x"05",  278 => x"15",  279 => x"00", 
         280 => x"93",  281 => x"85",  282 => x"15",  283 => x"00", 
         284 => x"63",  285 => x"14",  286 => x"d6",  287 => x"00", 
         288 => x"e3",  289 => x"16",  290 => x"06",  291 => x"fe", 
         292 => x"33",  293 => x"05",  294 => x"d6",  295 => x"40", 
         296 => x"67",  297 => x"80",  298 => x"00",  299 => x"00", 
         300 => x"13",  301 => x"01",  302 => x"01",  303 => x"ff", 
         304 => x"23",  305 => x"24",  306 => x"81",  307 => x"00", 
         308 => x"23",  309 => x"26",  310 => x"11",  311 => x"00", 
         312 => x"93",  313 => x"07",  314 => x"00",  315 => x"00", 
         316 => x"13",  317 => x"04",  318 => x"05",  319 => x"00", 
         320 => x"63",  321 => x"88",  322 => x"07",  323 => x"00", 
         324 => x"93",  325 => x"05",  326 => x"00",  327 => x"00", 
         328 => x"97",  329 => x"00",  330 => x"00",  331 => x"00", 
         332 => x"e7",  333 => x"00",  334 => x"00",  335 => x"00", 
         336 => x"03",  337 => x"25",  338 => x"80",  339 => x"28", 
         340 => x"83",  341 => x"27",  342 => x"85",  343 => x"02", 
         344 => x"63",  345 => x"84",  346 => x"07",  347 => x"00", 
         348 => x"e7",  349 => x"80",  350 => x"07",  351 => x"00", 
         352 => x"13",  353 => x"05",  354 => x"04",  355 => x"00", 
         356 => x"ef",  357 => x"00",  358 => x"80",  359 => x"0c", 
         360 => x"13",  361 => x"01",  362 => x"01",  363 => x"ff", 
         364 => x"23",  365 => x"24",  366 => x"81",  367 => x"00", 
         368 => x"23",  369 => x"22",  370 => x"91",  371 => x"00", 
         372 => x"93",  373 => x"07",  374 => x"c0",  375 => x"28", 
         376 => x"13",  377 => x"04",  378 => x"c0",  379 => x"28", 
         380 => x"33",  381 => x"04",  382 => x"f4",  383 => x"40", 
         384 => x"23",  385 => x"20",  386 => x"21",  387 => x"01", 
         388 => x"23",  389 => x"26",  390 => x"11",  391 => x"00", 
         392 => x"13",  393 => x"54",  394 => x"24",  395 => x"40", 
         396 => x"93",  397 => x"04",  398 => x"c0",  399 => x"28", 
         400 => x"13",  401 => x"09",  402 => x"00",  403 => x"00", 
         404 => x"63",  405 => x"1c",  406 => x"89",  407 => x"02", 
         408 => x"93",  409 => x"07",  410 => x"c0",  411 => x"28", 
         412 => x"13",  413 => x"04",  414 => x"c0",  415 => x"28", 
         416 => x"33",  417 => x"04",  418 => x"f4",  419 => x"40", 
         420 => x"13",  421 => x"54",  422 => x"24",  423 => x"40", 
         424 => x"93",  425 => x"04",  426 => x"c0",  427 => x"28", 
         428 => x"13",  429 => x"09",  430 => x"00",  431 => x"00", 
         432 => x"63",  433 => x"18",  434 => x"89",  435 => x"02", 
         436 => x"83",  437 => x"20",  438 => x"c1",  439 => x"00", 
         440 => x"03",  441 => x"24",  442 => x"81",  443 => x"00", 
         444 => x"83",  445 => x"24",  446 => x"41",  447 => x"00", 
         448 => x"03",  449 => x"29",  450 => x"01",  451 => x"00", 
         452 => x"13",  453 => x"01",  454 => x"01",  455 => x"01", 
         456 => x"67",  457 => x"80",  458 => x"00",  459 => x"00", 
         460 => x"83",  461 => x"a7",  462 => x"04",  463 => x"00", 
         464 => x"13",  465 => x"09",  466 => x"19",  467 => x"00", 
         468 => x"93",  469 => x"84",  470 => x"44",  471 => x"00", 
         472 => x"e7",  473 => x"80",  474 => x"07",  475 => x"00", 
         476 => x"6f",  477 => x"f0",  478 => x"9f",  479 => x"fb", 
         480 => x"83",  481 => x"a7",  482 => x"04",  483 => x"00", 
         484 => x"13",  485 => x"09",  486 => x"19",  487 => x"00", 
         488 => x"93",  489 => x"84",  490 => x"44",  491 => x"00", 
         492 => x"e7",  493 => x"80",  494 => x"07",  495 => x"00", 
         496 => x"6f",  497 => x"f0",  498 => x"1f",  499 => x"fc", 
         500 => x"93",  501 => x"07",  502 => x"05",  503 => x"00", 
         504 => x"03",  505 => x"c7",  506 => x"05",  507 => x"00", 
         508 => x"93",  509 => x"87",  510 => x"17",  511 => x"00", 
         512 => x"93",  513 => x"85",  514 => x"15",  515 => x"00", 
         516 => x"a3",  517 => x"8f",  518 => x"e7",  519 => x"fe", 
         520 => x"e3",  521 => x"18",  522 => x"07",  523 => x"fe", 
         524 => x"67",  525 => x"80",  526 => x"00",  527 => x"00", 
         528 => x"93",  529 => x"07",  530 => x"05",  531 => x"00", 
         532 => x"03",  533 => x"c7",  534 => x"07",  535 => x"00", 
         536 => x"93",  537 => x"87",  538 => x"17",  539 => x"00", 
         540 => x"e3",  541 => x"1c",  542 => x"07",  543 => x"fe", 
         544 => x"33",  545 => x"85",  546 => x"a7",  547 => x"40", 
         548 => x"13",  549 => x"05",  550 => x"f5",  551 => x"ff", 
         552 => x"67",  553 => x"80",  554 => x"00",  555 => x"00", 
         556 => x"93",  557 => x"08",  558 => x"d0",  559 => x"05", 
         560 => x"73",  561 => x"00",  562 => x"00",  563 => x"00", 
         564 => x"63",  565 => x"52",  566 => x"05",  567 => x"02", 
         568 => x"13",  569 => x"01",  570 => x"01",  571 => x"ff", 
         572 => x"23",  573 => x"24",  574 => x"81",  575 => x"00", 
         576 => x"13",  577 => x"04",  578 => x"05",  579 => x"00", 
         580 => x"23",  581 => x"26",  582 => x"11",  583 => x"00", 
         584 => x"33",  585 => x"04",  586 => x"80",  587 => x"40", 
         588 => x"ef",  589 => x"00",  590 => x"00",  591 => x"01", 
         592 => x"23",  593 => x"20",  594 => x"85",  595 => x"00", 
         596 => x"6f",  597 => x"00",  598 => x"00",  599 => x"00", 
         600 => x"6f",  601 => x"00",  602 => x"00",  603 => x"00", 
         604 => x"b7",  605 => x"07",  606 => x"00",  607 => x"20", 
         608 => x"03",  609 => x"a5",  610 => x"07",  611 => x"06", 
         612 => x"67",  613 => x"80",  614 => x"00",  615 => x"00", 
         616 => x"48",  617 => x"65",  618 => x"6c",  619 => x"6c", 
         620 => x"6f",  621 => x"00",  622 => x"00",  623 => x"00", 
         624 => x"48",  625 => x"65",  626 => x"6c",  627 => x"6c", 
         628 => x"6f",  629 => x"20",  630 => x"64",  631 => x"69", 
         632 => x"74",  633 => x"20",  634 => x"69",  635 => x"73", 
         636 => x"20",  637 => x"65",  638 => x"65",  639 => x"6e", 
         640 => x"20",  641 => x"73",  642 => x"74",  643 => x"72", 
         644 => x"69",  645 => x"6e",  646 => x"67",  647 => x"00", 
         648 => x"00",  649 => x"00",  650 => x"00",  651 => x"20", 
         652 => x"00",  653 => x"00",  654 => x"00",  655 => x"00", 
         656 => x"00",  657 => x"00",  658 => x"00",  659 => x"00", 
         660 => x"00",  661 => x"00",  662 => x"00",  663 => x"00", 
         664 => x"00",  665 => x"00",  666 => x"00",  667 => x"00", 
         668 => x"00",  669 => x"00",  670 => x"00",  671 => x"00", 
         672 => x"00",  673 => x"00",  674 => x"00",  675 => x"00", 
         676 => x"00",  677 => x"00",  678 => x"00",  679 => x"00", 
         680 => x"00",  681 => x"00",  682 => x"00",  683 => x"00", 
         684 => x"00",  685 => x"00",  686 => x"00",  687 => x"00", 
         688 => x"00",  689 => x"00",  690 => x"00",  691 => x"00", 
         692 => x"00",  693 => x"00",  694 => x"00",  695 => x"00", 
         696 => x"00",  697 => x"00",  698 => x"00",  699 => x"00", 
         700 => x"00",  701 => x"00",  702 => x"00",  703 => x"00", 
         704 => x"00",  705 => x"00",  706 => x"00",  707 => x"00", 
         708 => x"00",  709 => x"00",  710 => x"00",  711 => x"00", 
         712 => x"00",  713 => x"00",  714 => x"00",  715 => x"00", 
         716 => x"00",  717 => x"00",  718 => x"00",  719 => x"00", 
         720 => x"00",  721 => x"00",  722 => x"00",  723 => x"00", 
         724 => x"00",  725 => x"00",  726 => x"00",  727 => x"00", 
         728 => x"00",  729 => x"00",  730 => x"00",  731 => x"00", 
         732 => x"00",  733 => x"00",  734 => x"00",  735 => x"00", 
         736 => x"00",  737 => x"00",  738 => x"00",  739 => x"00", 
         740 => x"00",  741 => x"00",  742 => x"00",  743 => x"00", 
         744 => x"00",  745 => x"00",  746 => x"00",  747 => x"00", 
         748 => x"00",  749 => x"00",  750 => x"00",  751 => x"20", 
        others => (others => '-')
    );
end package processor_common_rom;
