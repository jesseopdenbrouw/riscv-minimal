-- srec2vhdl table generator
-- for input file main.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"93828206",
           6 => x"73905230",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef10803c",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"938505fe",
          21 => x"13050500",
          22 => x"ef100038",
          23 => x"ef10c06f",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10403e",
          29 => x"ef10406a",
          30 => x"6f000000",
          31 => x"37170000",
          32 => x"b70700f0",
          33 => x"13077745",
          34 => x"23a2e702",
          35 => x"13070004",
          36 => x"23a4e702",
          37 => x"67800000",
          38 => x"1375f50f",
          39 => x"b70700f0",
          40 => x"23a0a702",
          41 => x"370700f0",
          42 => x"8327c702",
          43 => x"93f70701",
          44 => x"e38c07fe",
          45 => x"67800000",
          46 => x"63060502",
          47 => x"83470500",
          48 => x"63820702",
          49 => x"370700f0",
          50 => x"13051500",
          51 => x"2320f702",
          52 => x"8327c702",
          53 => x"93f70701",
          54 => x"e38c07fe",
          55 => x"83470500",
          56 => x"e39407fe",
          57 => x"67800000",
          58 => x"370700f0",
          59 => x"8327c702",
          60 => x"93f74700",
          61 => x"e38c07fe",
          62 => x"03250702",
          63 => x"1375f50f",
          64 => x"67800000",
          65 => x"130101ff",
          66 => x"373e0000",
          67 => x"370700f0",
          68 => x"930e0500",
          69 => x"138ff5ff",
          70 => x"23268100",
          71 => x"13050000",
          72 => x"130e4ebe",
          73 => x"13070702",
          74 => x"13035001",
          75 => x"93027000",
          76 => x"930fe005",
          77 => x"9305f007",
          78 => x"93082000",
          79 => x"13082001",
          80 => x"b7330000",
          81 => x"1306f007",
          82 => x"8327c700",
          83 => x"93f74700",
          84 => x"e38c07fe",
          85 => x"03240700",
          86 => x"9376f40f",
          87 => x"636ed302",
          88 => x"63fed802",
          89 => x"9387d6ff",
          90 => x"636af802",
          91 => x"93972700",
          92 => x"b307fe00",
          93 => x"83a70700",
          94 => x"67800700",
          95 => x"1305f5ff",
          96 => x"6308050c",
          97 => x"2320c700",
          98 => x"8327c700",
          99 => x"93f70701",
         100 => x"e38c07fe",
         101 => x"6ff09ffe",
         102 => x"638cb606",
         103 => x"635ae50d",
         104 => x"1374f40f",
         105 => x"930704fe",
         106 => x"93f7f70f",
         107 => x"e3eefff8",
         108 => x"b387ae00",
         109 => x"23808700",
         110 => x"13051500",
         111 => x"2320d700",
         112 => x"8327c700",
         113 => x"93f70701",
         114 => x"e38c07fe",
         115 => x"6ff0dff7",
         116 => x"b38eae00",
         117 => x"b7360000",
         118 => x"23800e00",
         119 => x"9307d000",
         120 => x"938606e6",
         121 => x"370700f0",
         122 => x"93861600",
         123 => x"2320f702",
         124 => x"8327c702",
         125 => x"93f70701",
         126 => x"e38c07fe",
         127 => x"83c70600",
         128 => x"e39407fe",
         129 => x"0324c100",
         130 => x"13010101",
         131 => x"67800000",
         132 => x"63040504",
         133 => x"2320b700",
         134 => x"8327c700",
         135 => x"93f70701",
         136 => x"e38c07fe",
         137 => x"1305f5ff",
         138 => x"6ff01ff2",
         139 => x"9307c003",
         140 => x"938683f2",
         141 => x"93861600",
         142 => x"2320f700",
         143 => x"8327c700",
         144 => x"93f70701",
         145 => x"e38c07fe",
         146 => x"83c70600",
         147 => x"e39407fe",
         148 => x"13050000",
         149 => x"6ff05fef",
         150 => x"23205700",
         151 => x"8327c700",
         152 => x"93f70701",
         153 => x"e38c07fe",
         154 => x"13050000",
         155 => x"6ff0dfed",
         156 => x"23205700",
         157 => x"8327c700",
         158 => x"93f70701",
         159 => x"e38c07fe",
         160 => x"6ff09fec",
         161 => x"1375f50f",
         162 => x"b70700f0",
         163 => x"23a0a702",
         164 => x"370700f0",
         165 => x"8327c702",
         166 => x"93f70701",
         167 => x"e38c07fe",
         168 => x"13051000",
         169 => x"67800000",
         170 => x"370700f0",
         171 => x"8327c702",
         172 => x"93f74700",
         173 => x"e38c07fe",
         174 => x"03250702",
         175 => x"1375f50f",
         176 => x"67800000",
         177 => x"13050000",
         178 => x"67800000",
         179 => x"13050000",
         180 => x"67800000",
         181 => x"130101f8",
         182 => x"23221100",
         183 => x"23242100",
         184 => x"23263100",
         185 => x"23284100",
         186 => x"232a5100",
         187 => x"232c6100",
         188 => x"232e7100",
         189 => x"23208102",
         190 => x"23229102",
         191 => x"2324a102",
         192 => x"2326b102",
         193 => x"2328c102",
         194 => x"232ad102",
         195 => x"232ce102",
         196 => x"232ef102",
         197 => x"23200105",
         198 => x"23221105",
         199 => x"23242105",
         200 => x"23263105",
         201 => x"23284105",
         202 => x"232a5105",
         203 => x"232c6105",
         204 => x"232e7105",
         205 => x"23208107",
         206 => x"23229107",
         207 => x"2324a107",
         208 => x"2326b107",
         209 => x"2328c107",
         210 => x"232ad107",
         211 => x"232ce107",
         212 => x"232ef107",
         213 => x"f3272034",
         214 => x"37070080",
         215 => x"93067700",
         216 => x"6388d70c",
         217 => x"9306b000",
         218 => x"63e4f602",
         219 => x"13071000",
         220 => x"637cf70a",
         221 => x"63eaf60a",
         222 => x"37370000",
         223 => x"93972700",
         224 => x"130707c3",
         225 => x"b387e700",
         226 => x"83a70700",
         227 => x"67800700",
         228 => x"93061701",
         229 => x"6384d70a",
         230 => x"13072701",
         231 => x"6396e708",
         232 => x"ef008038",
         233 => x"03258102",
         234 => x"832fc107",
         235 => x"032f8107",
         236 => x"832e4107",
         237 => x"032e0107",
         238 => x"832dc106",
         239 => x"032d8106",
         240 => x"832c4106",
         241 => x"032c0106",
         242 => x"832bc105",
         243 => x"032b8105",
         244 => x"832a4105",
         245 => x"032a0105",
         246 => x"8329c104",
         247 => x"03298104",
         248 => x"83284104",
         249 => x"03280104",
         250 => x"8327c103",
         251 => x"03278103",
         252 => x"83264103",
         253 => x"03260103",
         254 => x"8325c102",
         255 => x"83244102",
         256 => x"03240102",
         257 => x"8323c101",
         258 => x"03238101",
         259 => x"83224101",
         260 => x"03220101",
         261 => x"8321c100",
         262 => x"03218100",
         263 => x"83204100",
         264 => x"13010108",
         265 => x"73002030",
         266 => x"03258102",
         267 => x"6ff0dff7",
         268 => x"ef00c02a",
         269 => x"03258102",
         270 => x"6ff01ff7",
         271 => x"ef00c026",
         272 => x"03258102",
         273 => x"6ff05ff6",
         274 => x"9307600d",
         275 => x"6388f814",
         276 => x"9307900a",
         277 => x"6382f818",
         278 => x"63cc1703",
         279 => x"938878fc",
         280 => x"93074002",
         281 => x"63e81705",
         282 => x"b7370000",
         283 => x"938707c6",
         284 => x"93982800",
         285 => x"b388f800",
         286 => x"83a70800",
         287 => x"67800700",
         288 => x"13050100",
         289 => x"ef00c01b",
         290 => x"03258102",
         291 => x"6ff0dff1",
         292 => x"938808c0",
         293 => x"9307f000",
         294 => x"63ee1701",
         295 => x"b7370000",
         296 => x"938747cf",
         297 => x"93982800",
         298 => x"b388f800",
         299 => x"83a70800",
         300 => x"67800700",
         301 => x"ef10c025",
         302 => x"93078005",
         303 => x"2320f500",
         304 => x"9307f0ff",
         305 => x"13850700",
         306 => x"6ff01fee",
         307 => x"b7270000",
         308 => x"23a2f500",
         309 => x"93070000",
         310 => x"13850700",
         311 => x"6ff0dfec",
         312 => x"93070000",
         313 => x"13850700",
         314 => x"6ff01fec",
         315 => x"ef104022",
         316 => x"93079000",
         317 => x"2320f500",
         318 => x"9307f0ff",
         319 => x"13850700",
         320 => x"6ff09fea",
         321 => x"ef10c020",
         322 => x"9307f001",
         323 => x"2320f500",
         324 => x"9307f0ff",
         325 => x"13850700",
         326 => x"6ff01fe9",
         327 => x"ef10401f",
         328 => x"9307d000",
         329 => x"2320f500",
         330 => x"9307f0ff",
         331 => x"13850700",
         332 => x"6ff09fe7",
         333 => x"ef10c01d",
         334 => x"93072000",
         335 => x"2320f500",
         336 => x"9307f0ff",
         337 => x"13850700",
         338 => x"6ff01fe6",
         339 => x"13090600",
         340 => x"13840500",
         341 => x"635cc000",
         342 => x"b384c500",
         343 => x"03450400",
         344 => x"13041400",
         345 => x"eff01fd2",
         346 => x"e39a84fe",
         347 => x"13050900",
         348 => x"6ff09fe3",
         349 => x"13090600",
         350 => x"13840500",
         351 => x"e358c0fe",
         352 => x"b384c500",
         353 => x"eff05fd2",
         354 => x"2300a400",
         355 => x"13041400",
         356 => x"e31a94fe",
         357 => x"13050900",
         358 => x"6ff01fe1",
         359 => x"63180500",
         360 => x"13858189",
         361 => x"13050500",
         362 => x"6ff01fe0",
         363 => x"b7870020",
         364 => x"93870700",
         365 => x"13070040",
         366 => x"b387e740",
         367 => x"e364f5fe",
         368 => x"ef100015",
         369 => x"9307c000",
         370 => x"2320f500",
         371 => x"1305f0ff",
         372 => x"13050500",
         373 => x"6ff05fdd",
         374 => x"13090000",
         375 => x"93040500",
         376 => x"13040900",
         377 => x"93090900",
         378 => x"93070900",
         379 => x"732410c8",
         380 => x"f32910c0",
         381 => x"f32710c8",
         382 => x"e31af4fe",
         383 => x"37460f00",
         384 => x"13060624",
         385 => x"93060000",
         386 => x"13850900",
         387 => x"93050400",
         388 => x"ef00501e",
         389 => x"37460f00",
         390 => x"23a4a400",
         391 => x"13060624",
         392 => x"93060000",
         393 => x"13850900",
         394 => x"93050400",
         395 => x"ef008059",
         396 => x"23a0a400",
         397 => x"23a2b400",
         398 => x"13050900",
         399 => x"6ff0dfd6",
         400 => x"37350000",
         401 => x"130101ff",
         402 => x"130545f3",
         403 => x"23261100",
         404 => x"23248100",
         405 => x"23229100",
         406 => x"23202101",
         407 => x"eff0dfa5",
         408 => x"73294034",
         409 => x"93040002",
         410 => x"37040080",
         411 => x"33758900",
         412 => x"3335a000",
         413 => x"13050503",
         414 => x"9384f4ff",
         415 => x"eff0dfa1",
         416 => x"13541400",
         417 => x"e39404fe",
         418 => x"03248100",
         419 => x"8320c100",
         420 => x"83244100",
         421 => x"03290100",
         422 => x"37350000",
         423 => x"130505e6",
         424 => x"13010101",
         425 => x"6ff05fa1",
         426 => x"b70700f0",
         427 => x"03a74708",
         428 => x"1377f7fe",
         429 => x"23a2e708",
         430 => x"03a74700",
         431 => x"13471700",
         432 => x"23a2e700",
         433 => x"67800000",
         434 => x"370700f0",
         435 => x"83274700",
         436 => x"93e70720",
         437 => x"2322f700",
         438 => x"6f000000",
         439 => x"b70700f0",
         440 => x"83a6470f",
         441 => x"03a6070f",
         442 => x"03a7470f",
         443 => x"e31ad7fe",
         444 => x"b7860100",
         445 => x"9305f0ff",
         446 => x"9386066a",
         447 => x"23aeb70e",
         448 => x"b306d600",
         449 => x"23acb70e",
         450 => x"33b6c600",
         451 => x"23acd70e",
         452 => x"3306e600",
         453 => x"23aec70e",
         454 => x"03a74700",
         455 => x"13472700",
         456 => x"23a2e700",
         457 => x"67800000",
         458 => x"370700f0",
         459 => x"8327c702",
         460 => x"93f74700",
         461 => x"638a0700",
         462 => x"83274700",
         463 => x"93c74700",
         464 => x"2322f700",
         465 => x"83270702",
         466 => x"67800000",
         467 => x"13030500",
         468 => x"138e0500",
         469 => x"93080000",
         470 => x"63dc0500",
         471 => x"b337a000",
         472 => x"330eb040",
         473 => x"330efe40",
         474 => x"3303a040",
         475 => x"9308f0ff",
         476 => x"63dc0600",
         477 => x"b337c000",
         478 => x"b306d040",
         479 => x"93c8f8ff",
         480 => x"b386f640",
         481 => x"3306c040",
         482 => x"13070600",
         483 => x"13080300",
         484 => x"93070e00",
         485 => x"639c0628",
         486 => x"b7350000",
         487 => x"938545d3",
         488 => x"6376ce0e",
         489 => x"b7060100",
         490 => x"6378d60c",
         491 => x"93360610",
         492 => x"93c61600",
         493 => x"93963600",
         494 => x"3355d600",
         495 => x"b385a500",
         496 => x"83c50500",
         497 => x"13050002",
         498 => x"b386d500",
         499 => x"b305d540",
         500 => x"630cd500",
         501 => x"b317be00",
         502 => x"b356d300",
         503 => x"3317b600",
         504 => x"b3e7f600",
         505 => x"3318b300",
         506 => x"93550701",
         507 => x"33deb702",
         508 => x"13160701",
         509 => x"13560601",
         510 => x"b3f7b702",
         511 => x"13050e00",
         512 => x"3303c603",
         513 => x"93960701",
         514 => x"93570801",
         515 => x"b3e7d700",
         516 => x"63fe6700",
         517 => x"b387e700",
         518 => x"1305feff",
         519 => x"63e8e700",
         520 => x"63f66700",
         521 => x"1305eeff",
         522 => x"b387e700",
         523 => x"b3876740",
         524 => x"33d3b702",
         525 => x"13180801",
         526 => x"13580801",
         527 => x"b3f7b702",
         528 => x"b3066602",
         529 => x"93970701",
         530 => x"3368f800",
         531 => x"93070300",
         532 => x"637cd800",
         533 => x"33080701",
         534 => x"9307f3ff",
         535 => x"6366e800",
         536 => x"6374d800",
         537 => x"9307e3ff",
         538 => x"13150501",
         539 => x"3365f500",
         540 => x"93050000",
         541 => x"6f00000e",
         542 => x"37050001",
         543 => x"93060001",
         544 => x"e36ca6f2",
         545 => x"93068001",
         546 => x"6ff01ff3",
         547 => x"63140600",
         548 => x"73001000",
         549 => x"b7070100",
         550 => x"637af60c",
         551 => x"93360610",
         552 => x"93c61600",
         553 => x"93963600",
         554 => x"b357d600",
         555 => x"b385f500",
         556 => x"83c70500",
         557 => x"b387d700",
         558 => x"93060002",
         559 => x"b385f640",
         560 => x"6390f60c",
         561 => x"b307ce40",
         562 => x"93051000",
         563 => x"13530701",
         564 => x"b3de6702",
         565 => x"13160701",
         566 => x"13560601",
         567 => x"93560801",
         568 => x"b3f76702",
         569 => x"13850e00",
         570 => x"330ed603",
         571 => x"93970701",
         572 => x"b3e7f600",
         573 => x"63fec701",
         574 => x"b387e700",
         575 => x"1385feff",
         576 => x"63e8e700",
         577 => x"63f6c701",
         578 => x"1385eeff",
         579 => x"b387e700",
         580 => x"b387c741",
         581 => x"33de6702",
         582 => x"13180801",
         583 => x"13580801",
         584 => x"b3f76702",
         585 => x"b306c603",
         586 => x"93970701",
         587 => x"3368f800",
         588 => x"93070e00",
         589 => x"637cd800",
         590 => x"33080701",
         591 => x"9307feff",
         592 => x"6366e800",
         593 => x"6374d800",
         594 => x"9307eeff",
         595 => x"13150501",
         596 => x"3365f500",
         597 => x"638a0800",
         598 => x"b337a000",
         599 => x"b305b040",
         600 => x"b385f540",
         601 => x"3305a040",
         602 => x"67800000",
         603 => x"b7070001",
         604 => x"93060001",
         605 => x"e36af6f2",
         606 => x"93068001",
         607 => x"6ff0dff2",
         608 => x"3317b600",
         609 => x"b356fe00",
         610 => x"13550701",
         611 => x"331ebe00",
         612 => x"b357f300",
         613 => x"b3e7c701",
         614 => x"33dea602",
         615 => x"13160701",
         616 => x"13560601",
         617 => x"3318b300",
         618 => x"b3f6a602",
         619 => x"3303c603",
         620 => x"93950601",
         621 => x"93d60701",
         622 => x"b3e6b600",
         623 => x"93050e00",
         624 => x"63fe6600",
         625 => x"b386e600",
         626 => x"9305feff",
         627 => x"63e8e600",
         628 => x"63f66600",
         629 => x"9305eeff",
         630 => x"b386e600",
         631 => x"b3866640",
         632 => x"33d3a602",
         633 => x"93970701",
         634 => x"93d70701",
         635 => x"b3f6a602",
         636 => x"33066602",
         637 => x"93960601",
         638 => x"b3e7d700",
         639 => x"93060300",
         640 => x"63fec700",
         641 => x"b387e700",
         642 => x"9306f3ff",
         643 => x"63e8e700",
         644 => x"63f6c700",
         645 => x"9306e3ff",
         646 => x"b387e700",
         647 => x"93950501",
         648 => x"b387c740",
         649 => x"b3e5d500",
         650 => x"6ff05fea",
         651 => x"6366de18",
         652 => x"b7070100",
         653 => x"63f4f604",
         654 => x"13b70610",
         655 => x"13471700",
         656 => x"13173700",
         657 => x"b7370000",
         658 => x"b3d5e600",
         659 => x"938747d3",
         660 => x"b387b700",
         661 => x"83c70700",
         662 => x"b387e700",
         663 => x"13070002",
         664 => x"b305f740",
         665 => x"6316f702",
         666 => x"13051000",
         667 => x"e3e4c6ef",
         668 => x"3335c300",
         669 => x"13451500",
         670 => x"6ff0dfed",
         671 => x"b7070001",
         672 => x"13070001",
         673 => x"e3e0f6fc",
         674 => x"13078001",
         675 => x"6ff09ffb",
         676 => x"3357f600",
         677 => x"b396b600",
         678 => x"b366d700",
         679 => x"3357fe00",
         680 => x"331ebe00",
         681 => x"b357f300",
         682 => x"b3e7c701",
         683 => x"13de0601",
         684 => x"335fc703",
         685 => x"13980601",
         686 => x"13580801",
         687 => x"3316b600",
         688 => x"3377c703",
         689 => x"b30ee803",
         690 => x"13150701",
         691 => x"13d70701",
         692 => x"3367a700",
         693 => x"13050f00",
         694 => x"637ed701",
         695 => x"3307d700",
         696 => x"1305ffff",
         697 => x"6368d700",
         698 => x"6376d701",
         699 => x"1305efff",
         700 => x"3307d700",
         701 => x"3307d741",
         702 => x"b35ec703",
         703 => x"93970701",
         704 => x"93d70701",
         705 => x"3377c703",
         706 => x"3308d803",
         707 => x"13170701",
         708 => x"b3e7e700",
         709 => x"13870e00",
         710 => x"63fe0701",
         711 => x"b387d700",
         712 => x"1387feff",
         713 => x"63e8d700",
         714 => x"63f60701",
         715 => x"1387eeff",
         716 => x"b387d700",
         717 => x"13150501",
         718 => x"b70e0100",
         719 => x"3365e500",
         720 => x"9386feff",
         721 => x"3377d500",
         722 => x"b3870741",
         723 => x"b376d600",
         724 => x"13580501",
         725 => x"13560601",
         726 => x"330ed702",
         727 => x"b306d802",
         728 => x"3307c702",
         729 => x"3308c802",
         730 => x"3306d700",
         731 => x"13570e01",
         732 => x"3307c700",
         733 => x"6374d700",
         734 => x"3308d801",
         735 => x"93560701",
         736 => x"b3860601",
         737 => x"63e6d702",
         738 => x"e394d7ce",
         739 => x"b7070100",
         740 => x"9387f7ff",
         741 => x"3377f700",
         742 => x"13170701",
         743 => x"337efe00",
         744 => x"3313b300",
         745 => x"3307c701",
         746 => x"93050000",
         747 => x"e374e3da",
         748 => x"1305f5ff",
         749 => x"6ff0dfcb",
         750 => x"93050000",
         751 => x"13050000",
         752 => x"6ff05fd9",
         753 => x"13030500",
         754 => x"93880500",
         755 => x"13070600",
         756 => x"13080500",
         757 => x"93870500",
         758 => x"63920628",
         759 => x"b7350000",
         760 => x"938545d3",
         761 => x"63f6c80e",
         762 => x"b7060100",
         763 => x"6378d60c",
         764 => x"93360610",
         765 => x"93c61600",
         766 => x"93963600",
         767 => x"3355d600",
         768 => x"b385a500",
         769 => x"83c50500",
         770 => x"13050002",
         771 => x"b386d500",
         772 => x"b305d540",
         773 => x"630cd500",
         774 => x"b397b800",
         775 => x"b356d300",
         776 => x"3317b600",
         777 => x"b3e7f600",
         778 => x"3318b300",
         779 => x"93550701",
         780 => x"33d3b702",
         781 => x"13160701",
         782 => x"13560601",
         783 => x"b3f7b702",
         784 => x"13050300",
         785 => x"b3086602",
         786 => x"93960701",
         787 => x"93570801",
         788 => x"b3e7d700",
         789 => x"63fe1701",
         790 => x"b387e700",
         791 => x"1305f3ff",
         792 => x"63e8e700",
         793 => x"63f61701",
         794 => x"1305e3ff",
         795 => x"b387e700",
         796 => x"b3871741",
         797 => x"b3d8b702",
         798 => x"13180801",
         799 => x"13580801",
         800 => x"b3f7b702",
         801 => x"b3061603",
         802 => x"93970701",
         803 => x"3368f800",
         804 => x"93870800",
         805 => x"637cd800",
         806 => x"33080701",
         807 => x"9387f8ff",
         808 => x"6366e800",
         809 => x"6374d800",
         810 => x"9387e8ff",
         811 => x"13150501",
         812 => x"3365f500",
         813 => x"93050000",
         814 => x"67800000",
         815 => x"37050001",
         816 => x"93060001",
         817 => x"e36ca6f2",
         818 => x"93068001",
         819 => x"6ff01ff3",
         820 => x"63140600",
         821 => x"73001000",
         822 => x"b7070100",
         823 => x"6370f60c",
         824 => x"93360610",
         825 => x"93c61600",
         826 => x"93963600",
         827 => x"b357d600",
         828 => x"b385f500",
         829 => x"83c70500",
         830 => x"b387d700",
         831 => x"93060002",
         832 => x"b385f640",
         833 => x"6396f60a",
         834 => x"b387c840",
         835 => x"93051000",
         836 => x"93580701",
         837 => x"33de1703",
         838 => x"13160701",
         839 => x"13560601",
         840 => x"93560801",
         841 => x"b3f71703",
         842 => x"13050e00",
         843 => x"3303c603",
         844 => x"93970701",
         845 => x"b3e7f600",
         846 => x"63fe6700",
         847 => x"b387e700",
         848 => x"1305feff",
         849 => x"63e8e700",
         850 => x"63f66700",
         851 => x"1305eeff",
         852 => x"b387e700",
         853 => x"b3876740",
         854 => x"33d31703",
         855 => x"13180801",
         856 => x"13580801",
         857 => x"b3f71703",
         858 => x"b3066602",
         859 => x"93970701",
         860 => x"3368f800",
         861 => x"93070300",
         862 => x"637cd800",
         863 => x"33080701",
         864 => x"9307f3ff",
         865 => x"6366e800",
         866 => x"6374d800",
         867 => x"9307e3ff",
         868 => x"13150501",
         869 => x"3365f500",
         870 => x"67800000",
         871 => x"b7070001",
         872 => x"93060001",
         873 => x"e364f6f4",
         874 => x"93068001",
         875 => x"6ff01ff4",
         876 => x"3317b600",
         877 => x"b3d6f800",
         878 => x"13550701",
         879 => x"b357f300",
         880 => x"3318b300",
         881 => x"33d3a602",
         882 => x"13160701",
         883 => x"b398b800",
         884 => x"13560601",
         885 => x"b3e71701",
         886 => x"b3f6a602",
         887 => x"b3086602",
         888 => x"93950601",
         889 => x"93d60701",
         890 => x"b3e6b600",
         891 => x"93050300",
         892 => x"63fe1601",
         893 => x"b386e600",
         894 => x"9305f3ff",
         895 => x"63e8e600",
         896 => x"63f61601",
         897 => x"9305e3ff",
         898 => x"b386e600",
         899 => x"b3861641",
         900 => x"b3d8a602",
         901 => x"93970701",
         902 => x"93d70701",
         903 => x"b3f6a602",
         904 => x"33061603",
         905 => x"93960601",
         906 => x"b3e7d700",
         907 => x"93860800",
         908 => x"63fec700",
         909 => x"b387e700",
         910 => x"9386f8ff",
         911 => x"63e8e700",
         912 => x"63f6c700",
         913 => x"9386e8ff",
         914 => x"b387e700",
         915 => x"93950501",
         916 => x"b387c740",
         917 => x"b3e5d500",
         918 => x"6ff09feb",
         919 => x"63e6d518",
         920 => x"b7070100",
         921 => x"63f4f604",
         922 => x"13b70610",
         923 => x"13471700",
         924 => x"13173700",
         925 => x"b7370000",
         926 => x"b3d5e600",
         927 => x"938747d3",
         928 => x"b387b700",
         929 => x"83c70700",
         930 => x"b387e700",
         931 => x"13070002",
         932 => x"b305f740",
         933 => x"6316f702",
         934 => x"13051000",
         935 => x"e3ee16e1",
         936 => x"3335c300",
         937 => x"13451500",
         938 => x"67800000",
         939 => x"b7070001",
         940 => x"13070001",
         941 => x"e3e0f6fc",
         942 => x"13078001",
         943 => x"6ff09ffb",
         944 => x"3357f600",
         945 => x"b396b600",
         946 => x"b366d700",
         947 => x"33d7f800",
         948 => x"b398b800",
         949 => x"b357f300",
         950 => x"b3e71701",
         951 => x"93d80601",
         952 => x"b35e1703",
         953 => x"13980601",
         954 => x"13580801",
         955 => x"3316b600",
         956 => x"33771703",
         957 => x"330ed803",
         958 => x"13150701",
         959 => x"13d70701",
         960 => x"3367a700",
         961 => x"13850e00",
         962 => x"637ec701",
         963 => x"3307d700",
         964 => x"1385feff",
         965 => x"6368d700",
         966 => x"6376c701",
         967 => x"1385eeff",
         968 => x"3307d700",
         969 => x"3307c741",
         970 => x"335e1703",
         971 => x"93970701",
         972 => x"93d70701",
         973 => x"33771703",
         974 => x"3308c803",
         975 => x"13170701",
         976 => x"b3e7e700",
         977 => x"13070e00",
         978 => x"63fe0701",
         979 => x"b387d700",
         980 => x"1307feff",
         981 => x"63e8d700",
         982 => x"63f60701",
         983 => x"1307eeff",
         984 => x"b387d700",
         985 => x"13150501",
         986 => x"370e0100",
         987 => x"3365e500",
         988 => x"9306feff",
         989 => x"3377d500",
         990 => x"b3870741",
         991 => x"b376d600",
         992 => x"13580501",
         993 => x"13560601",
         994 => x"b308d702",
         995 => x"b306d802",
         996 => x"3307c702",
         997 => x"3308c802",
         998 => x"3306d700",
         999 => x"13d70801",
        1000 => x"3307c700",
        1001 => x"6374d700",
        1002 => x"3308c801",
        1003 => x"93560701",
        1004 => x"b3860601",
        1005 => x"63e6d702",
        1006 => x"e39ed7ce",
        1007 => x"b7070100",
        1008 => x"9387f7ff",
        1009 => x"3377f700",
        1010 => x"13170701",
        1011 => x"b3f8f800",
        1012 => x"3313b300",
        1013 => x"33071701",
        1014 => x"93050000",
        1015 => x"e37ee3cc",
        1016 => x"1305f5ff",
        1017 => x"6ff01fcd",
        1018 => x"93050000",
        1019 => x"13050000",
        1020 => x"67800000",
        1021 => x"13080600",
        1022 => x"93070500",
        1023 => x"13870500",
        1024 => x"63960620",
        1025 => x"b7380000",
        1026 => x"938848d3",
        1027 => x"63fcc50c",
        1028 => x"b7060100",
        1029 => x"637ed60a",
        1030 => x"93360610",
        1031 => x"93c61600",
        1032 => x"93963600",
        1033 => x"3353d600",
        1034 => x"b3886800",
        1035 => x"83c80800",
        1036 => x"13030002",
        1037 => x"b386d800",
        1038 => x"b308d340",
        1039 => x"630cd300",
        1040 => x"33971501",
        1041 => x"b356d500",
        1042 => x"33181601",
        1043 => x"33e7e600",
        1044 => x"b3171501",
        1045 => x"13560801",
        1046 => x"b356c702",
        1047 => x"13150801",
        1048 => x"13550501",
        1049 => x"3377c702",
        1050 => x"b386a602",
        1051 => x"93150701",
        1052 => x"13d70701",
        1053 => x"3367b700",
        1054 => x"637ad700",
        1055 => x"33070701",
        1056 => x"63660701",
        1057 => x"6374d700",
        1058 => x"33070701",
        1059 => x"3307d740",
        1060 => x"b356c702",
        1061 => x"3377c702",
        1062 => x"b386a602",
        1063 => x"93970701",
        1064 => x"13170701",
        1065 => x"93d70701",
        1066 => x"b3e7e700",
        1067 => x"63fad700",
        1068 => x"b3870701",
        1069 => x"63e60701",
        1070 => x"63f4d700",
        1071 => x"b3870701",
        1072 => x"b387d740",
        1073 => x"33d51701",
        1074 => x"93050000",
        1075 => x"67800000",
        1076 => x"37030001",
        1077 => x"93060001",
        1078 => x"e36666f4",
        1079 => x"93068001",
        1080 => x"6ff05ff4",
        1081 => x"63140600",
        1082 => x"73001000",
        1083 => x"37070100",
        1084 => x"637ee606",
        1085 => x"93360610",
        1086 => x"93c61600",
        1087 => x"93963600",
        1088 => x"3357d600",
        1089 => x"b388e800",
        1090 => x"03c70800",
        1091 => x"3307d700",
        1092 => x"93060002",
        1093 => x"b388e640",
        1094 => x"6394e606",
        1095 => x"3387c540",
        1096 => x"93550801",
        1097 => x"3356b702",
        1098 => x"13150801",
        1099 => x"13550501",
        1100 => x"93d60701",
        1101 => x"3377b702",
        1102 => x"3306a602",
        1103 => x"13170701",
        1104 => x"33e7e600",
        1105 => x"637ac700",
        1106 => x"33070701",
        1107 => x"63660701",
        1108 => x"6374c700",
        1109 => x"33070701",
        1110 => x"3307c740",
        1111 => x"b356b702",
        1112 => x"3377b702",
        1113 => x"b386a602",
        1114 => x"6ff05ff3",
        1115 => x"37070001",
        1116 => x"93060001",
        1117 => x"e366e6f8",
        1118 => x"93068001",
        1119 => x"6ff05ff8",
        1120 => x"33181601",
        1121 => x"b3d6e500",
        1122 => x"b3171501",
        1123 => x"b3951501",
        1124 => x"3357e500",
        1125 => x"13550801",
        1126 => x"3367b700",
        1127 => x"b3d5a602",
        1128 => x"13130801",
        1129 => x"13530301",
        1130 => x"b3f6a602",
        1131 => x"b3856502",
        1132 => x"13960601",
        1133 => x"93560701",
        1134 => x"b3e6c600",
        1135 => x"63fab600",
        1136 => x"b3860601",
        1137 => x"63e60601",
        1138 => x"63f4b600",
        1139 => x"b3860601",
        1140 => x"b386b640",
        1141 => x"33d6a602",
        1142 => x"13170701",
        1143 => x"13570701",
        1144 => x"b3f6a602",
        1145 => x"33066602",
        1146 => x"93960601",
        1147 => x"3367d700",
        1148 => x"637ac700",
        1149 => x"33070701",
        1150 => x"63660701",
        1151 => x"6374c700",
        1152 => x"33070701",
        1153 => x"3307c740",
        1154 => x"6ff09ff1",
        1155 => x"63e4d51c",
        1156 => x"37080100",
        1157 => x"63fe0605",
        1158 => x"13b80610",
        1159 => x"13481800",
        1160 => x"13183800",
        1161 => x"b7380000",
        1162 => x"33d30601",
        1163 => x"938848d3",
        1164 => x"b3886800",
        1165 => x"83c80800",
        1166 => x"13030002",
        1167 => x"b3880801",
        1168 => x"33081341",
        1169 => x"63101305",
        1170 => x"63e4b600",
        1171 => x"636cc500",
        1172 => x"3306c540",
        1173 => x"b386d540",
        1174 => x"3337c500",
        1175 => x"3387e640",
        1176 => x"93070600",
        1177 => x"13850700",
        1178 => x"93050700",
        1179 => x"67800000",
        1180 => x"b7080001",
        1181 => x"13080001",
        1182 => x"e3e616fb",
        1183 => x"13088001",
        1184 => x"6ff05ffa",
        1185 => x"b3960601",
        1186 => x"33531601",
        1187 => x"3363d300",
        1188 => x"135e0301",
        1189 => x"b3d61501",
        1190 => x"33dfc603",
        1191 => x"13170301",
        1192 => x"13570701",
        1193 => x"b3970501",
        1194 => x"b3551501",
        1195 => x"b3e5f500",
        1196 => x"93d70501",
        1197 => x"33160601",
        1198 => x"33150501",
        1199 => x"b3f6c603",
        1200 => x"b30ee703",
        1201 => x"93960601",
        1202 => x"b3e7d700",
        1203 => x"93060f00",
        1204 => x"63fed701",
        1205 => x"b3876700",
        1206 => x"9306ffff",
        1207 => x"63e86700",
        1208 => x"63f6d701",
        1209 => x"9306efff",
        1210 => x"b3876700",
        1211 => x"b387d741",
        1212 => x"b3dec703",
        1213 => x"93950501",
        1214 => x"93d50501",
        1215 => x"b3f7c703",
        1216 => x"3307d703",
        1217 => x"93970701",
        1218 => x"b3e5f500",
        1219 => x"93870e00",
        1220 => x"63fee500",
        1221 => x"b3856500",
        1222 => x"9387feff",
        1223 => x"63e86500",
        1224 => x"63f6e500",
        1225 => x"9387eeff",
        1226 => x"b3856500",
        1227 => x"93960601",
        1228 => x"370f0100",
        1229 => x"b3e6f600",
        1230 => x"9307ffff",
        1231 => x"135e0601",
        1232 => x"b385e540",
        1233 => x"33f7f600",
        1234 => x"93d60601",
        1235 => x"b377f600",
        1236 => x"b30ef702",
        1237 => x"b387f602",
        1238 => x"3307c703",
        1239 => x"b386c603",
        1240 => x"330ef700",
        1241 => x"13d70e01",
        1242 => x"3307c701",
        1243 => x"6374f700",
        1244 => x"b386e601",
        1245 => x"93570701",
        1246 => x"b387d700",
        1247 => x"b7060100",
        1248 => x"9386f6ff",
        1249 => x"3377d700",
        1250 => x"13170701",
        1251 => x"b3fede00",
        1252 => x"3307d701",
        1253 => x"63e6f500",
        1254 => x"639ef500",
        1255 => x"637ce500",
        1256 => x"3306c740",
        1257 => x"3337c700",
        1258 => x"33076700",
        1259 => x"b387e740",
        1260 => x"13070600",
        1261 => x"3307e540",
        1262 => x"3335e500",
        1263 => x"b385f540",
        1264 => x"b385a540",
        1265 => x"b3981501",
        1266 => x"33570701",
        1267 => x"33e5e800",
        1268 => x"b3d50501",
        1269 => x"67800000",
        1270 => x"13030500",
        1271 => x"630e0600",
        1272 => x"83830500",
        1273 => x"23007300",
        1274 => x"1306f6ff",
        1275 => x"13031300",
        1276 => x"93851500",
        1277 => x"e31606fe",
        1278 => x"67800000",
        1279 => x"13030500",
        1280 => x"630a0600",
        1281 => x"2300b300",
        1282 => x"1306f6ff",
        1283 => x"13031300",
        1284 => x"e31a06fe",
        1285 => x"67800000",
        1286 => x"630c0602",
        1287 => x"13030500",
        1288 => x"93061000",
        1289 => x"636ab500",
        1290 => x"9306f0ff",
        1291 => x"1307f6ff",
        1292 => x"3303e300",
        1293 => x"b385e500",
        1294 => x"83830500",
        1295 => x"23007300",
        1296 => x"1306f6ff",
        1297 => x"3303d300",
        1298 => x"b385d500",
        1299 => x"e31606fe",
        1300 => x"67800000",
        1301 => x"130101f8",
        1302 => x"232c8106",
        1303 => x"23263107",
        1304 => x"232e1106",
        1305 => x"232a9106",
        1306 => x"23282107",
        1307 => x"23244107",
        1308 => x"23225107",
        1309 => x"23206107",
        1310 => x"232e7105",
        1311 => x"232c8105",
        1312 => x"232a9105",
        1313 => x"2328a105",
        1314 => x"2326b105",
        1315 => x"93090500",
        1316 => x"13840500",
        1317 => x"232c0100",
        1318 => x"232e0100",
        1319 => x"23200102",
        1320 => x"23220102",
        1321 => x"23240102",
        1322 => x"23260102",
        1323 => x"23280102",
        1324 => x"232a0102",
        1325 => x"232c0102",
        1326 => x"232e0102",
        1327 => x"97f2ffff",
        1328 => x"938282e1",
        1329 => x"73905230",
        1330 => x"efe05fbb",
        1331 => x"b7877d01",
        1332 => x"370700f0",
        1333 => x"9387f783",
        1334 => x"2326f708",
        1335 => x"93071001",
        1336 => x"2320f708",
        1337 => x"93020008",
        1338 => x"73904230",
        1339 => x"b7220000",
        1340 => x"93828280",
        1341 => x"73900230",
        1342 => x"37390000",
        1343 => x"130509e6",
        1344 => x"efe09fbb",
        1345 => x"63543003",
        1346 => x"9384f9ff",
        1347 => x"9309f0ff",
        1348 => x"03250400",
        1349 => x"9384f4ff",
        1350 => x"13044400",
        1351 => x"efe0dfb9",
        1352 => x"130509e6",
        1353 => x"efe05fb9",
        1354 => x"e39434ff",
        1355 => x"37350000",
        1356 => x"b7faeeee",
        1357 => x"130545e3",
        1358 => x"b7040010",
        1359 => x"37190000",
        1360 => x"1384faee",
        1361 => x"efe05fb7",
        1362 => x"130c0000",
        1363 => x"b73b0000",
        1364 => x"9384f4ff",
        1365 => x"130bf000",
        1366 => x"938aeaee",
        1367 => x"130909e1",
        1368 => x"93090000",
        1369 => x"130a0019",
        1370 => x"93050000",
        1371 => x"13058100",
        1372 => x"ef008035",
        1373 => x"130c1c00",
        1374 => x"63020502",
        1375 => x"e3164cff",
        1376 => x"73001000",
        1377 => x"93050000",
        1378 => x"13058100",
        1379 => x"130c0000",
        1380 => x"ef008033",
        1381 => x"130c1c00",
        1382 => x"e31205fe",
        1383 => x"832c8100",
        1384 => x"8325c100",
        1385 => x"13060900",
        1386 => x"93d7cc01",
        1387 => x"13974500",
        1388 => x"b367f700",
        1389 => x"b3f79700",
        1390 => x"33f79c00",
        1391 => x"13d5f541",
        1392 => x"13d88501",
        1393 => x"3307f700",
        1394 => x"33070701",
        1395 => x"9377d500",
        1396 => x"3307f700",
        1397 => x"33776703",
        1398 => x"937725ff",
        1399 => x"93860900",
        1400 => x"13850c00",
        1401 => x"3307f700",
        1402 => x"b387ec40",
        1403 => x"1357f741",
        1404 => x"33b8fc00",
        1405 => x"3387e540",
        1406 => x"33070741",
        1407 => x"b3885703",
        1408 => x"33078702",
        1409 => x"33b88702",
        1410 => x"33071701",
        1411 => x"b3878702",
        1412 => x"33070701",
        1413 => x"1358f741",
        1414 => x"13783800",
        1415 => x"b307f800",
        1416 => x"33b80701",
        1417 => x"3307e800",
        1418 => x"1318e701",
        1419 => x"93d72700",
        1420 => x"b367f800",
        1421 => x"93582740",
        1422 => x"13984800",
        1423 => x"13d3c701",
        1424 => x"33636800",
        1425 => x"33739300",
        1426 => x"33f89700",
        1427 => x"13de8801",
        1428 => x"1357f741",
        1429 => x"33086800",
        1430 => x"3308c801",
        1431 => x"1373d700",
        1432 => x"33086800",
        1433 => x"33786803",
        1434 => x"137727ff",
        1435 => x"139d4700",
        1436 => x"330dfd40",
        1437 => x"131d2d00",
        1438 => x"338dac41",
        1439 => x"3308e800",
        1440 => x"33870741",
        1441 => x"1358f841",
        1442 => x"33b3e700",
        1443 => x"b3880841",
        1444 => x"b3886840",
        1445 => x"b3888802",
        1446 => x"33035703",
        1447 => x"33388702",
        1448 => x"b3886800",
        1449 => x"33078702",
        1450 => x"b3880801",
        1451 => x"13d8f841",
        1452 => x"13783800",
        1453 => x"3307e800",
        1454 => x"33380701",
        1455 => x"33081801",
        1456 => x"1318e801",
        1457 => x"13572700",
        1458 => x"3367e800",
        1459 => x"13184700",
        1460 => x"3307e840",
        1461 => x"13172700",
        1462 => x"b38de740",
        1463 => x"eff00f87",
        1464 => x"83260101",
        1465 => x"13070500",
        1466 => x"13080d00",
        1467 => x"93870d00",
        1468 => x"13860c00",
        1469 => x"93854be6",
        1470 => x"13058101",
        1471 => x"ef00c015",
        1472 => x"13058101",
        1473 => x"efe05f9b",
        1474 => x"e3104ce7",
        1475 => x"6ff05fe7",
        1476 => x"03a5c187",
        1477 => x"67800000",
        1478 => x"130101ff",
        1479 => x"23248100",
        1480 => x"23261100",
        1481 => x"93070000",
        1482 => x"13040500",
        1483 => x"63880700",
        1484 => x"93050000",
        1485 => x"97000000",
        1486 => x"e7000000",
        1487 => x"b7370000",
        1488 => x"03a5c7fd",
        1489 => x"83278502",
        1490 => x"63840700",
        1491 => x"e7800700",
        1492 => x"13050400",
        1493 => x"ef108033",
        1494 => x"130101ff",
        1495 => x"23248100",
        1496 => x"23229100",
        1497 => x"37340000",
        1498 => x"b7340000",
        1499 => x"938704fe",
        1500 => x"130404fe",
        1501 => x"3304f440",
        1502 => x"23202101",
        1503 => x"23261100",
        1504 => x"13542440",
        1505 => x"938404fe",
        1506 => x"13090000",
        1507 => x"63108904",
        1508 => x"b7340000",
        1509 => x"37340000",
        1510 => x"938704fe",
        1511 => x"130404fe",
        1512 => x"3304f440",
        1513 => x"13542440",
        1514 => x"938404fe",
        1515 => x"13090000",
        1516 => x"63188902",
        1517 => x"8320c100",
        1518 => x"03248100",
        1519 => x"83244100",
        1520 => x"03290100",
        1521 => x"13010101",
        1522 => x"67800000",
        1523 => x"83a70400",
        1524 => x"13091900",
        1525 => x"93844400",
        1526 => x"e7800700",
        1527 => x"6ff01ffb",
        1528 => x"83a70400",
        1529 => x"13091900",
        1530 => x"93844400",
        1531 => x"e7800700",
        1532 => x"6ff01ffc",
        1533 => x"130101f6",
        1534 => x"232af108",
        1535 => x"b7070080",
        1536 => x"93c7f7ff",
        1537 => x"232ef100",
        1538 => x"2328f100",
        1539 => x"b707ffff",
        1540 => x"2326d108",
        1541 => x"2324b100",
        1542 => x"232cb100",
        1543 => x"93878720",
        1544 => x"9306c108",
        1545 => x"93058100",
        1546 => x"232e1106",
        1547 => x"232af100",
        1548 => x"2328e108",
        1549 => x"232c0109",
        1550 => x"232e1109",
        1551 => x"2322d100",
        1552 => x"ef004041",
        1553 => x"83278100",
        1554 => x"23800700",
        1555 => x"8320c107",
        1556 => x"1301010a",
        1557 => x"67800000",
        1558 => x"130101f6",
        1559 => x"232af108",
        1560 => x"b7070080",
        1561 => x"93c7f7ff",
        1562 => x"232ef100",
        1563 => x"2328f100",
        1564 => x"b707ffff",
        1565 => x"93878720",
        1566 => x"232af100",
        1567 => x"2324a100",
        1568 => x"232ca100",
        1569 => x"03a5c187",
        1570 => x"2324c108",
        1571 => x"2326d108",
        1572 => x"13860500",
        1573 => x"93068108",
        1574 => x"93058100",
        1575 => x"232e1106",
        1576 => x"2328e108",
        1577 => x"232c0109",
        1578 => x"232e1109",
        1579 => x"2322d100",
        1580 => x"ef00403a",
        1581 => x"83278100",
        1582 => x"23800700",
        1583 => x"8320c107",
        1584 => x"1301010a",
        1585 => x"67800000",
        1586 => x"13860500",
        1587 => x"93050500",
        1588 => x"03a5c187",
        1589 => x"6f004000",
        1590 => x"130101ff",
        1591 => x"23248100",
        1592 => x"23229100",
        1593 => x"13040500",
        1594 => x"13850500",
        1595 => x"93050600",
        1596 => x"23261100",
        1597 => x"23a20188",
        1598 => x"ef10401c",
        1599 => x"9307f0ff",
        1600 => x"6318f500",
        1601 => x"83a74188",
        1602 => x"63840700",
        1603 => x"2320f400",
        1604 => x"8320c100",
        1605 => x"03248100",
        1606 => x"83244100",
        1607 => x"13010101",
        1608 => x"67800000",
        1609 => x"130101fe",
        1610 => x"23282101",
        1611 => x"03a98500",
        1612 => x"232c8100",
        1613 => x"23263101",
        1614 => x"23244101",
        1615 => x"23225101",
        1616 => x"232e1100",
        1617 => x"232a9100",
        1618 => x"23206101",
        1619 => x"83aa0500",
        1620 => x"13840500",
        1621 => x"130a0600",
        1622 => x"93890600",
        1623 => x"63ec2609",
        1624 => x"83d7c500",
        1625 => x"13f70748",
        1626 => x"63040708",
        1627 => x"03274401",
        1628 => x"93043000",
        1629 => x"83a50501",
        1630 => x"b384e402",
        1631 => x"13072000",
        1632 => x"b38aba40",
        1633 => x"130b0500",
        1634 => x"b3c4e402",
        1635 => x"13871600",
        1636 => x"33075701",
        1637 => x"63f4e400",
        1638 => x"93040700",
        1639 => x"93f70740",
        1640 => x"6386070a",
        1641 => x"93850400",
        1642 => x"13050b00",
        1643 => x"ef001065",
        1644 => x"13090500",
        1645 => x"630c050a",
        1646 => x"83250401",
        1647 => x"13860a00",
        1648 => x"eff09fa1",
        1649 => x"8357c400",
        1650 => x"93f7f7b7",
        1651 => x"93e70708",
        1652 => x"2316f400",
        1653 => x"23282401",
        1654 => x"232a9400",
        1655 => x"33095901",
        1656 => x"b3845441",
        1657 => x"23202401",
        1658 => x"23249400",
        1659 => x"13890900",
        1660 => x"63f42901",
        1661 => x"13890900",
        1662 => x"03250400",
        1663 => x"13060900",
        1664 => x"93050a00",
        1665 => x"eff05fa1",
        1666 => x"83278400",
        1667 => x"13050000",
        1668 => x"b3872741",
        1669 => x"2324f400",
        1670 => x"83270400",
        1671 => x"b3872701",
        1672 => x"2320f400",
        1673 => x"8320c101",
        1674 => x"03248101",
        1675 => x"83244101",
        1676 => x"03290101",
        1677 => x"8329c100",
        1678 => x"032a8100",
        1679 => x"832a4100",
        1680 => x"032b0100",
        1681 => x"13010102",
        1682 => x"67800000",
        1683 => x"13860400",
        1684 => x"13050b00",
        1685 => x"ef00906f",
        1686 => x"13090500",
        1687 => x"e31c05f6",
        1688 => x"83250401",
        1689 => x"13050b00",
        1690 => x"ef00d049",
        1691 => x"9307c000",
        1692 => x"2320fb00",
        1693 => x"8357c400",
        1694 => x"1305f0ff",
        1695 => x"93e70704",
        1696 => x"2316f400",
        1697 => x"6ff01ffa",
        1698 => x"83278600",
        1699 => x"130101fd",
        1700 => x"232e3101",
        1701 => x"23286101",
        1702 => x"23261102",
        1703 => x"23248102",
        1704 => x"23229102",
        1705 => x"23202103",
        1706 => x"232c4101",
        1707 => x"232a5101",
        1708 => x"23267101",
        1709 => x"23248101",
        1710 => x"23229101",
        1711 => x"2320a101",
        1712 => x"032b0600",
        1713 => x"93090600",
        1714 => x"63980712",
        1715 => x"13050000",
        1716 => x"8320c102",
        1717 => x"03248102",
        1718 => x"23a20900",
        1719 => x"83244102",
        1720 => x"03290102",
        1721 => x"8329c101",
        1722 => x"032a8101",
        1723 => x"832a4101",
        1724 => x"032b0101",
        1725 => x"832bc100",
        1726 => x"032c8100",
        1727 => x"832c4100",
        1728 => x"032d0100",
        1729 => x"13010103",
        1730 => x"67800000",
        1731 => x"832a0b00",
        1732 => x"032d4b00",
        1733 => x"130b8b00",
        1734 => x"03298400",
        1735 => x"832c0400",
        1736 => x"e3060dfe",
        1737 => x"63642d09",
        1738 => x"8357c400",
        1739 => x"13f70748",
        1740 => x"630e0706",
        1741 => x"83244401",
        1742 => x"83250401",
        1743 => x"b3849b02",
        1744 => x"b38cbc40",
        1745 => x"13871c00",
        1746 => x"3307a701",
        1747 => x"b3c48403",
        1748 => x"63f4e400",
        1749 => x"93040700",
        1750 => x"93f70740",
        1751 => x"638c070a",
        1752 => x"93850400",
        1753 => x"13050a00",
        1754 => x"ef005049",
        1755 => x"13090500",
        1756 => x"6302050c",
        1757 => x"83250401",
        1758 => x"13860c00",
        1759 => x"eff0df85",
        1760 => x"8357c400",
        1761 => x"93f7f7b7",
        1762 => x"93e70708",
        1763 => x"2316f400",
        1764 => x"23282401",
        1765 => x"232a9400",
        1766 => x"33099901",
        1767 => x"b3849441",
        1768 => x"23202401",
        1769 => x"23249400",
        1770 => x"13090d00",
        1771 => x"63742d01",
        1772 => x"13090d00",
        1773 => x"03250400",
        1774 => x"93850a00",
        1775 => x"13060900",
        1776 => x"eff09f85",
        1777 => x"83278400",
        1778 => x"b38aaa01",
        1779 => x"b3872741",
        1780 => x"2324f400",
        1781 => x"83270400",
        1782 => x"b3872701",
        1783 => x"2320f400",
        1784 => x"83a78900",
        1785 => x"b387a741",
        1786 => x"23a4f900",
        1787 => x"e38007ee",
        1788 => x"130d0000",
        1789 => x"6ff05ff2",
        1790 => x"130a0500",
        1791 => x"13840500",
        1792 => x"930a0000",
        1793 => x"130d0000",
        1794 => x"930b3000",
        1795 => x"130c2000",
        1796 => x"6ff09ff0",
        1797 => x"13860400",
        1798 => x"13050a00",
        1799 => x"ef001053",
        1800 => x"13090500",
        1801 => x"e31605f6",
        1802 => x"83250401",
        1803 => x"13050a00",
        1804 => x"ef00502d",
        1805 => x"9307c000",
        1806 => x"2320fa00",
        1807 => x"8357c400",
        1808 => x"1305f0ff",
        1809 => x"93e70704",
        1810 => x"2316f400",
        1811 => x"23a40900",
        1812 => x"6ff01fe8",
        1813 => x"83d7c500",
        1814 => x"130101f5",
        1815 => x"2324810a",
        1816 => x"2322910a",
        1817 => x"2320210b",
        1818 => x"232c4109",
        1819 => x"2326110a",
        1820 => x"232e3109",
        1821 => x"232a5109",
        1822 => x"23286109",
        1823 => x"23267109",
        1824 => x"23248109",
        1825 => x"23229109",
        1826 => x"2320a109",
        1827 => x"232eb107",
        1828 => x"93f70708",
        1829 => x"130a0500",
        1830 => x"13890500",
        1831 => x"93040600",
        1832 => x"13840600",
        1833 => x"63880706",
        1834 => x"83a70501",
        1835 => x"63940706",
        1836 => x"93050004",
        1837 => x"ef009034",
        1838 => x"2320a900",
        1839 => x"2328a900",
        1840 => x"63160504",
        1841 => x"9307c000",
        1842 => x"2320fa00",
        1843 => x"1305f0ff",
        1844 => x"8320c10a",
        1845 => x"0324810a",
        1846 => x"8324410a",
        1847 => x"0329010a",
        1848 => x"8329c109",
        1849 => x"032a8109",
        1850 => x"832a4109",
        1851 => x"032b0109",
        1852 => x"832bc108",
        1853 => x"032c8108",
        1854 => x"832c4108",
        1855 => x"032d0108",
        1856 => x"832dc107",
        1857 => x"1301010b",
        1858 => x"67800000",
        1859 => x"93070004",
        1860 => x"232af900",
        1861 => x"93070002",
        1862 => x"a304f102",
        1863 => x"93070003",
        1864 => x"23220102",
        1865 => x"2305f102",
        1866 => x"23268100",
        1867 => x"930c5002",
        1868 => x"373b0000",
        1869 => x"b73b0000",
        1870 => x"373d0000",
        1871 => x"372c0000",
        1872 => x"930a0000",
        1873 => x"13840400",
        1874 => x"83470400",
        1875 => x"63840700",
        1876 => x"639c970d",
        1877 => x"b30d9440",
        1878 => x"63069402",
        1879 => x"93860d00",
        1880 => x"13860400",
        1881 => x"93050900",
        1882 => x"13050a00",
        1883 => x"eff09fbb",
        1884 => x"9307f0ff",
        1885 => x"6306f524",
        1886 => x"83274102",
        1887 => x"b387b701",
        1888 => x"2322f102",
        1889 => x"83470400",
        1890 => x"638c0722",
        1891 => x"9307f0ff",
        1892 => x"93041400",
        1893 => x"23280100",
        1894 => x"232e0100",
        1895 => x"232af100",
        1896 => x"232c0100",
        1897 => x"a3090104",
        1898 => x"23240106",
        1899 => x"930d1000",
        1900 => x"83c50400",
        1901 => x"13065000",
        1902 => x"13058bf4",
        1903 => x"ef005012",
        1904 => x"83270101",
        1905 => x"13841400",
        1906 => x"63140506",
        1907 => x"13f70701",
        1908 => x"63060700",
        1909 => x"13070002",
        1910 => x"a309e104",
        1911 => x"13f78700",
        1912 => x"63060700",
        1913 => x"1307b002",
        1914 => x"a309e104",
        1915 => x"83c60400",
        1916 => x"1307a002",
        1917 => x"638ce604",
        1918 => x"8327c101",
        1919 => x"13840400",
        1920 => x"93060000",
        1921 => x"13069000",
        1922 => x"1305a000",
        1923 => x"03470400",
        1924 => x"93051400",
        1925 => x"130707fd",
        1926 => x"637ce608",
        1927 => x"63840604",
        1928 => x"232ef100",
        1929 => x"6f000004",
        1930 => x"13041400",
        1931 => x"6ff0dff1",
        1932 => x"13078bf4",
        1933 => x"3305e540",
        1934 => x"3395ad00",
        1935 => x"b3e7a700",
        1936 => x"2328f100",
        1937 => x"93040400",
        1938 => x"6ff09ff6",
        1939 => x"0327c100",
        1940 => x"93064700",
        1941 => x"03270700",
        1942 => x"2326d100",
        1943 => x"63400704",
        1944 => x"232ee100",
        1945 => x"03470400",
        1946 => x"9307e002",
        1947 => x"6316f708",
        1948 => x"03471400",
        1949 => x"9307a002",
        1950 => x"631af704",
        1951 => x"8327c100",
        1952 => x"13042400",
        1953 => x"13874700",
        1954 => x"83a70700",
        1955 => x"2326e100",
        1956 => x"63ca0702",
        1957 => x"232af100",
        1958 => x"6f000006",
        1959 => x"3307e040",
        1960 => x"93e72700",
        1961 => x"232ee100",
        1962 => x"2328f100",
        1963 => x"6ff09ffb",
        1964 => x"b387a702",
        1965 => x"13840500",
        1966 => x"93061000",
        1967 => x"b387e700",
        1968 => x"6ff0dff4",
        1969 => x"9307f0ff",
        1970 => x"6ff0dffc",
        1971 => x"13041400",
        1972 => x"232a0100",
        1973 => x"93060000",
        1974 => x"93070000",
        1975 => x"13069000",
        1976 => x"1305a000",
        1977 => x"03470400",
        1978 => x"93051400",
        1979 => x"130707fd",
        1980 => x"6372e608",
        1981 => x"e39006fa",
        1982 => x"83450400",
        1983 => x"13063000",
        1984 => x"13850bf5",
        1985 => x"ef00c07d",
        1986 => x"63020502",
        1987 => x"93870bf5",
        1988 => x"3305f540",
        1989 => x"83270101",
        1990 => x"13070004",
        1991 => x"3317a700",
        1992 => x"b3e7e700",
        1993 => x"13041400",
        1994 => x"2328f100",
        1995 => x"83450400",
        1996 => x"13066000",
        1997 => x"13054df5",
        1998 => x"93041400",
        1999 => x"2304b102",
        2000 => x"ef00007a",
        2001 => x"630a0508",
        2002 => x"63980a04",
        2003 => x"03270101",
        2004 => x"8327c100",
        2005 => x"13770710",
        2006 => x"63080702",
        2007 => x"93874700",
        2008 => x"2326f100",
        2009 => x"83274102",
        2010 => x"b3873701",
        2011 => x"2322f102",
        2012 => x"6ff05fdd",
        2013 => x"b387a702",
        2014 => x"13840500",
        2015 => x"93061000",
        2016 => x"b387e700",
        2017 => x"6ff01ff6",
        2018 => x"93877700",
        2019 => x"93f787ff",
        2020 => x"93878700",
        2021 => x"6ff0dffc",
        2022 => x"1307c100",
        2023 => x"93064c92",
        2024 => x"13060900",
        2025 => x"93050101",
        2026 => x"13050a00",
        2027 => x"97000000",
        2028 => x"e7000000",
        2029 => x"9307f0ff",
        2030 => x"93090500",
        2031 => x"e314f5fa",
        2032 => x"8357c900",
        2033 => x"1305f0ff",
        2034 => x"93f70704",
        2035 => x"e39207d0",
        2036 => x"03254102",
        2037 => x"6ff0dfcf",
        2038 => x"1307c100",
        2039 => x"93064c92",
        2040 => x"13060900",
        2041 => x"93050101",
        2042 => x"13050a00",
        2043 => x"ef00801b",
        2044 => x"6ff05ffc",
        2045 => x"130101fd",
        2046 => x"232c4101",
        2047 => x"83a70501",
        2048 => x"130a0700",
        2049 => x"03a78500",
        2050 => x"23248102",
        2051 => x"23202103",
        2052 => x"232e3101",
        2053 => x"232a5101",
        2054 => x"23261102",
        2055 => x"23229102",
        2056 => x"23286101",
        2057 => x"23267101",
        2058 => x"93090500",
        2059 => x"13840500",
        2060 => x"13090600",
        2061 => x"938a0600",
        2062 => x"63d4e700",
        2063 => x"93070700",
        2064 => x"2320f900",
        2065 => x"03473404",
        2066 => x"63060700",
        2067 => x"93871700",
        2068 => x"2320f900",
        2069 => x"83270400",
        2070 => x"93f70702",
        2071 => x"63880700",
        2072 => x"83270900",
        2073 => x"93872700",
        2074 => x"2320f900",
        2075 => x"83240400",
        2076 => x"93f46400",
        2077 => x"639e0400",
        2078 => x"130b9401",
        2079 => x"930bf0ff",
        2080 => x"8327c400",
        2081 => x"03270900",
        2082 => x"b387e740",
        2083 => x"63c2f408",
        2084 => x"83473404",
        2085 => x"b336f000",
        2086 => x"83270400",
        2087 => x"93f70702",
        2088 => x"6390070c",
        2089 => x"13063404",
        2090 => x"93850a00",
        2091 => x"13850900",
        2092 => x"e7000a00",
        2093 => x"9307f0ff",
        2094 => x"6308f506",
        2095 => x"83270400",
        2096 => x"13074000",
        2097 => x"93040000",
        2098 => x"93f76700",
        2099 => x"639ce700",
        2100 => x"8324c400",
        2101 => x"83270900",
        2102 => x"b384f440",
        2103 => x"63d40400",
        2104 => x"93040000",
        2105 => x"83278400",
        2106 => x"03270401",
        2107 => x"6356f700",
        2108 => x"b387e740",
        2109 => x"b384f400",
        2110 => x"13090000",
        2111 => x"1304a401",
        2112 => x"130bf0ff",
        2113 => x"63902409",
        2114 => x"13050000",
        2115 => x"6f000002",
        2116 => x"93061000",
        2117 => x"13060b00",
        2118 => x"93850a00",
        2119 => x"13850900",
        2120 => x"e7000a00",
        2121 => x"631a7503",
        2122 => x"1305f0ff",
        2123 => x"8320c102",
        2124 => x"03248102",
        2125 => x"83244102",
        2126 => x"03290102",
        2127 => x"8329c101",
        2128 => x"032a8101",
        2129 => x"832a4101",
        2130 => x"032b0101",
        2131 => x"832bc100",
        2132 => x"13010103",
        2133 => x"67800000",
        2134 => x"93841400",
        2135 => x"6ff05ff2",
        2136 => x"3307d400",
        2137 => x"13060003",
        2138 => x"a301c704",
        2139 => x"03475404",
        2140 => x"93871600",
        2141 => x"b307f400",
        2142 => x"93862600",
        2143 => x"a381e704",
        2144 => x"6ff05ff2",
        2145 => x"93061000",
        2146 => x"13060400",
        2147 => x"93850a00",
        2148 => x"13850900",
        2149 => x"e7000a00",
        2150 => x"e30865f9",
        2151 => x"13091900",
        2152 => x"6ff05ff6",
        2153 => x"130101fd",
        2154 => x"23248102",
        2155 => x"23229102",
        2156 => x"23202103",
        2157 => x"232e3101",
        2158 => x"23261102",
        2159 => x"232c4101",
        2160 => x"232a5101",
        2161 => x"23286101",
        2162 => x"83c88501",
        2163 => x"93078007",
        2164 => x"93040500",
        2165 => x"13840500",
        2166 => x"13090600",
        2167 => x"93890600",
        2168 => x"63ee1701",
        2169 => x"93072006",
        2170 => x"93863504",
        2171 => x"63ee1701",
        2172 => x"63840828",
        2173 => x"93078005",
        2174 => x"6388f822",
        2175 => x"930a2404",
        2176 => x"23011405",
        2177 => x"6f004004",
        2178 => x"9387d8f9",
        2179 => x"93f7f70f",
        2180 => x"13065001",
        2181 => x"e364f6fe",
        2182 => x"37360000",
        2183 => x"93972700",
        2184 => x"130646f8",
        2185 => x"b387c700",
        2186 => x"83a70700",
        2187 => x"67800700",
        2188 => x"83270700",
        2189 => x"938a2504",
        2190 => x"93864700",
        2191 => x"83a70700",
        2192 => x"2320d700",
        2193 => x"2381f504",
        2194 => x"93071000",
        2195 => x"6f008026",
        2196 => x"83a70500",
        2197 => x"03250700",
        2198 => x"13f60708",
        2199 => x"93054500",
        2200 => x"63060602",
        2201 => x"83270500",
        2202 => x"2320b700",
        2203 => x"37380000",
        2204 => x"63d80700",
        2205 => x"1307d002",
        2206 => x"b307f040",
        2207 => x"a301e404",
        2208 => x"1308c8f5",
        2209 => x"1307a000",
        2210 => x"6f008006",
        2211 => x"13f60704",
        2212 => x"83270500",
        2213 => x"2320b700",
        2214 => x"e30a06fc",
        2215 => x"93970701",
        2216 => x"93d70741",
        2217 => x"6ff09ffc",
        2218 => x"03a60500",
        2219 => x"83270700",
        2220 => x"13750608",
        2221 => x"93854700",
        2222 => x"63080500",
        2223 => x"2320b700",
        2224 => x"83a70700",
        2225 => x"6f004001",
        2226 => x"13760604",
        2227 => x"2320b700",
        2228 => x"e30806fe",
        2229 => x"83d70700",
        2230 => x"37380000",
        2231 => x"1307f006",
        2232 => x"1308c8f5",
        2233 => x"6388e814",
        2234 => x"1307a000",
        2235 => x"a3010404",
        2236 => x"03264400",
        2237 => x"2324c400",
        2238 => x"63480600",
        2239 => x"83250400",
        2240 => x"93f5b5ff",
        2241 => x"2320b400",
        2242 => x"63960700",
        2243 => x"938a0600",
        2244 => x"63040602",
        2245 => x"938a0600",
        2246 => x"33f6e702",
        2247 => x"938afaff",
        2248 => x"3306c800",
        2249 => x"03460600",
        2250 => x"2380ca00",
        2251 => x"13860700",
        2252 => x"b3d7e702",
        2253 => x"e372e6fe",
        2254 => x"93078000",
        2255 => x"6314f702",
        2256 => x"83270400",
        2257 => x"93f71700",
        2258 => x"638e0700",
        2259 => x"03274400",
        2260 => x"83270401",
        2261 => x"63c8e700",
        2262 => x"93070003",
        2263 => x"a38ffafe",
        2264 => x"938afaff",
        2265 => x"b3865641",
        2266 => x"2328d400",
        2267 => x"13870900",
        2268 => x"93060900",
        2269 => x"1306c100",
        2270 => x"93050400",
        2271 => x"13850400",
        2272 => x"eff05fc7",
        2273 => x"130af0ff",
        2274 => x"631c4513",
        2275 => x"1305f0ff",
        2276 => x"8320c102",
        2277 => x"03248102",
        2278 => x"83244102",
        2279 => x"03290102",
        2280 => x"8329c101",
        2281 => x"032a8101",
        2282 => x"832a4101",
        2283 => x"032b0101",
        2284 => x"13010103",
        2285 => x"67800000",
        2286 => x"83a70500",
        2287 => x"93e70702",
        2288 => x"23a0f500",
        2289 => x"37380000",
        2290 => x"93088007",
        2291 => x"130808f7",
        2292 => x"a3021405",
        2293 => x"03260400",
        2294 => x"83250700",
        2295 => x"13750608",
        2296 => x"83a70500",
        2297 => x"93854500",
        2298 => x"631a0500",
        2299 => x"13750604",
        2300 => x"63060500",
        2301 => x"93970701",
        2302 => x"93d70701",
        2303 => x"2320b700",
        2304 => x"13771600",
        2305 => x"63060700",
        2306 => x"13660602",
        2307 => x"2320c400",
        2308 => x"13070001",
        2309 => x"e39c07ec",
        2310 => x"03260400",
        2311 => x"1376f6fd",
        2312 => x"2320c400",
        2313 => x"6ff09fec",
        2314 => x"37380000",
        2315 => x"1308c8f5",
        2316 => x"6ff01ffa",
        2317 => x"13078000",
        2318 => x"6ff05feb",
        2319 => x"03a60500",
        2320 => x"83270700",
        2321 => x"83a54501",
        2322 => x"13780608",
        2323 => x"13854700",
        2324 => x"630a0800",
        2325 => x"2320a700",
        2326 => x"83a70700",
        2327 => x"23a0b700",
        2328 => x"6f008001",
        2329 => x"2320a700",
        2330 => x"13760604",
        2331 => x"83a70700",
        2332 => x"e30606fe",
        2333 => x"2390b700",
        2334 => x"23280400",
        2335 => x"938a0600",
        2336 => x"6ff0dfee",
        2337 => x"83270700",
        2338 => x"03a64500",
        2339 => x"93050000",
        2340 => x"93864700",
        2341 => x"2320d700",
        2342 => x"83aa0700",
        2343 => x"13850a00",
        2344 => x"ef000024",
        2345 => x"63060500",
        2346 => x"33055541",
        2347 => x"2322a400",
        2348 => x"83274400",
        2349 => x"2328f400",
        2350 => x"a3010404",
        2351 => x"6ff01feb",
        2352 => x"83260401",
        2353 => x"13860a00",
        2354 => x"93050900",
        2355 => x"13850400",
        2356 => x"e7800900",
        2357 => x"e30c45eb",
        2358 => x"83270400",
        2359 => x"93f72700",
        2360 => x"63940704",
        2361 => x"8327c100",
        2362 => x"0325c400",
        2363 => x"e352f5ea",
        2364 => x"13850700",
        2365 => x"6ff0dfe9",
        2366 => x"93061000",
        2367 => x"13860a00",
        2368 => x"93050900",
        2369 => x"13850400",
        2370 => x"e7800900",
        2371 => x"e30065e9",
        2372 => x"130a1a00",
        2373 => x"8327c400",
        2374 => x"0327c100",
        2375 => x"b387e740",
        2376 => x"e34cfafc",
        2377 => x"6ff01ffc",
        2378 => x"130a0000",
        2379 => x"930a9401",
        2380 => x"130bf0ff",
        2381 => x"6ff01ffe",
        2382 => x"130101ff",
        2383 => x"23248100",
        2384 => x"13840500",
        2385 => x"83a50500",
        2386 => x"23229100",
        2387 => x"23261100",
        2388 => x"93040500",
        2389 => x"63840500",
        2390 => x"eff01ffe",
        2391 => x"93050400",
        2392 => x"03248100",
        2393 => x"8320c100",
        2394 => x"13850400",
        2395 => x"83244100",
        2396 => x"13010101",
        2397 => x"6f000019",
        2398 => x"83a7c187",
        2399 => x"6380a716",
        2400 => x"83274502",
        2401 => x"130101fe",
        2402 => x"232c8100",
        2403 => x"232e1100",
        2404 => x"232a9100",
        2405 => x"23282101",
        2406 => x"23263101",
        2407 => x"13040500",
        2408 => x"63840702",
        2409 => x"83a7c700",
        2410 => x"93040000",
        2411 => x"13090008",
        2412 => x"6392070e",
        2413 => x"83274402",
        2414 => x"83a50700",
        2415 => x"63860500",
        2416 => x"13050400",
        2417 => x"ef000014",
        2418 => x"83254401",
        2419 => x"63860500",
        2420 => x"13050400",
        2421 => x"ef000013",
        2422 => x"83254402",
        2423 => x"63860500",
        2424 => x"13050400",
        2425 => x"ef000012",
        2426 => x"83258403",
        2427 => x"63860500",
        2428 => x"13050400",
        2429 => x"ef000011",
        2430 => x"8325c403",
        2431 => x"63860500",
        2432 => x"13050400",
        2433 => x"ef000010",
        2434 => x"83250404",
        2435 => x"63860500",
        2436 => x"13050400",
        2437 => x"ef00000f",
        2438 => x"8325c405",
        2439 => x"63860500",
        2440 => x"13050400",
        2441 => x"ef00000e",
        2442 => x"83258405",
        2443 => x"63860500",
        2444 => x"13050400",
        2445 => x"ef00000d",
        2446 => x"83254403",
        2447 => x"63860500",
        2448 => x"13050400",
        2449 => x"ef00000c",
        2450 => x"83278401",
        2451 => x"638a0706",
        2452 => x"83278402",
        2453 => x"13050400",
        2454 => x"e7800700",
        2455 => x"83258404",
        2456 => x"63800506",
        2457 => x"13050400",
        2458 => x"03248101",
        2459 => x"8320c101",
        2460 => x"83244101",
        2461 => x"03290101",
        2462 => x"8329c100",
        2463 => x"13010102",
        2464 => x"6ff09feb",
        2465 => x"b3859500",
        2466 => x"83a50500",
        2467 => x"63900502",
        2468 => x"93844400",
        2469 => x"83274402",
        2470 => x"83a5c700",
        2471 => x"e39424ff",
        2472 => x"13050400",
        2473 => x"ef000006",
        2474 => x"6ff0dff0",
        2475 => x"83a90500",
        2476 => x"13050400",
        2477 => x"ef000005",
        2478 => x"93850900",
        2479 => x"6ff01ffd",
        2480 => x"8320c101",
        2481 => x"03248101",
        2482 => x"83244101",
        2483 => x"03290101",
        2484 => x"8329c100",
        2485 => x"13010102",
        2486 => x"67800000",
        2487 => x"67800000",
        2488 => x"93f5f50f",
        2489 => x"3306c500",
        2490 => x"6316c500",
        2491 => x"13050000",
        2492 => x"67800000",
        2493 => x"83470500",
        2494 => x"e38cb7fe",
        2495 => x"13051500",
        2496 => x"6ff09ffe",
        2497 => x"638a050e",
        2498 => x"83a7c5ff",
        2499 => x"130101fe",
        2500 => x"232c8100",
        2501 => x"232e1100",
        2502 => x"1384c5ff",
        2503 => x"63d40700",
        2504 => x"3304f400",
        2505 => x"2326a100",
        2506 => x"ef000034",
        2507 => x"83a78188",
        2508 => x"0325c100",
        2509 => x"639e0700",
        2510 => x"23220400",
        2511 => x"23a48188",
        2512 => x"03248101",
        2513 => x"8320c101",
        2514 => x"13010102",
        2515 => x"6f000032",
        2516 => x"6374f402",
        2517 => x"03260400",
        2518 => x"b306c400",
        2519 => x"639ad700",
        2520 => x"83a60700",
        2521 => x"83a74700",
        2522 => x"b386c600",
        2523 => x"2320d400",
        2524 => x"2322f400",
        2525 => x"6ff09ffc",
        2526 => x"13870700",
        2527 => x"83a74700",
        2528 => x"63840700",
        2529 => x"e37af4fe",
        2530 => x"83260700",
        2531 => x"3306d700",
        2532 => x"63188602",
        2533 => x"03260400",
        2534 => x"b386c600",
        2535 => x"2320d700",
        2536 => x"3306d700",
        2537 => x"e39ec7f8",
        2538 => x"03a60700",
        2539 => x"83a74700",
        2540 => x"b306d600",
        2541 => x"2320d700",
        2542 => x"2322f700",
        2543 => x"6ff05ff8",
        2544 => x"6378c400",
        2545 => x"9307c000",
        2546 => x"2320f500",
        2547 => x"6ff05ff7",
        2548 => x"03260400",
        2549 => x"b306c400",
        2550 => x"639ad700",
        2551 => x"83a60700",
        2552 => x"83a74700",
        2553 => x"b386c600",
        2554 => x"2320d400",
        2555 => x"2322f400",
        2556 => x"23228700",
        2557 => x"6ff0dff4",
        2558 => x"67800000",
        2559 => x"130101fe",
        2560 => x"232a9100",
        2561 => x"93843500",
        2562 => x"93f4c4ff",
        2563 => x"23282101",
        2564 => x"232e1100",
        2565 => x"232c8100",
        2566 => x"23263101",
        2567 => x"93848400",
        2568 => x"9307c000",
        2569 => x"13090500",
        2570 => x"63f4f406",
        2571 => x"9304c000",
        2572 => x"63e2b406",
        2573 => x"13050900",
        2574 => x"ef000023",
        2575 => x"03a78188",
        2576 => x"93868188",
        2577 => x"13040700",
        2578 => x"631a0406",
        2579 => x"1384c188",
        2580 => x"83270400",
        2581 => x"639a0700",
        2582 => x"93050000",
        2583 => x"13050900",
        2584 => x"ef00001c",
        2585 => x"2320a400",
        2586 => x"93850400",
        2587 => x"13050900",
        2588 => x"ef00001b",
        2589 => x"9309f0ff",
        2590 => x"631a350b",
        2591 => x"9307c000",
        2592 => x"2320f900",
        2593 => x"13050900",
        2594 => x"ef00401e",
        2595 => x"6f000001",
        2596 => x"e3d004fa",
        2597 => x"9307c000",
        2598 => x"2320f900",
        2599 => x"13050000",
        2600 => x"8320c101",
        2601 => x"03248101",
        2602 => x"83244101",
        2603 => x"03290101",
        2604 => x"8329c100",
        2605 => x"13010102",
        2606 => x"67800000",
        2607 => x"83270400",
        2608 => x"b3879740",
        2609 => x"63ce0704",
        2610 => x"1306b000",
        2611 => x"637af600",
        2612 => x"2320f400",
        2613 => x"3304f400",
        2614 => x"23209400",
        2615 => x"6f000001",
        2616 => x"83274400",
        2617 => x"631a8702",
        2618 => x"23a0f600",
        2619 => x"13050900",
        2620 => x"ef00c017",
        2621 => x"1305b400",
        2622 => x"93074400",
        2623 => x"137585ff",
        2624 => x"3307f540",
        2625 => x"e30ef5f8",
        2626 => x"3304e400",
        2627 => x"b387a740",
        2628 => x"2320f400",
        2629 => x"6ff0dff8",
        2630 => x"2322f700",
        2631 => x"6ff01ffd",
        2632 => x"13070400",
        2633 => x"03244400",
        2634 => x"6ff01ff2",
        2635 => x"13043500",
        2636 => x"1374c4ff",
        2637 => x"e30285fa",
        2638 => x"b305a440",
        2639 => x"13050900",
        2640 => x"ef00000e",
        2641 => x"e31a35f9",
        2642 => x"6ff05ff3",
        2643 => x"130101fe",
        2644 => x"232c8100",
        2645 => x"232e1100",
        2646 => x"232a9100",
        2647 => x"23282101",
        2648 => x"23263101",
        2649 => x"23244101",
        2650 => x"13040600",
        2651 => x"63940502",
        2652 => x"03248101",
        2653 => x"8320c101",
        2654 => x"83244101",
        2655 => x"03290101",
        2656 => x"8329c100",
        2657 => x"032a8100",
        2658 => x"93050600",
        2659 => x"13010102",
        2660 => x"6ff0dfe6",
        2661 => x"63180602",
        2662 => x"eff0dfd6",
        2663 => x"93040000",
        2664 => x"8320c101",
        2665 => x"03248101",
        2666 => x"03290101",
        2667 => x"8329c100",
        2668 => x"032a8100",
        2669 => x"13850400",
        2670 => x"83244101",
        2671 => x"13010102",
        2672 => x"67800000",
        2673 => x"130a0500",
        2674 => x"13890500",
        2675 => x"ef00400a",
        2676 => x"93090500",
        2677 => x"63688500",
        2678 => x"93571500",
        2679 => x"93040900",
        2680 => x"e3e087fc",
        2681 => x"93050400",
        2682 => x"13050a00",
        2683 => x"eff01fe1",
        2684 => x"93040500",
        2685 => x"e30605fa",
        2686 => x"13060400",
        2687 => x"63f48900",
        2688 => x"13860900",
        2689 => x"93050900",
        2690 => x"13850400",
        2691 => x"efe0df9c",
        2692 => x"93050900",
        2693 => x"13050a00",
        2694 => x"eff0dfce",
        2695 => x"6ff05ff8",
        2696 => x"130101ff",
        2697 => x"23248100",
        2698 => x"23229100",
        2699 => x"13040500",
        2700 => x"13850500",
        2701 => x"23261100",
        2702 => x"23a20188",
        2703 => x"ef00000c",
        2704 => x"9307f0ff",
        2705 => x"6318f500",
        2706 => x"83a74188",
        2707 => x"63840700",
        2708 => x"2320f400",
        2709 => x"8320c100",
        2710 => x"03248100",
        2711 => x"83244100",
        2712 => x"13010101",
        2713 => x"67800000",
        2714 => x"67800000",
        2715 => x"67800000",
        2716 => x"83a7c5ff",
        2717 => x"1385c7ff",
        2718 => x"63d80700",
        2719 => x"b385a500",
        2720 => x"83a70500",
        2721 => x"3305f500",
        2722 => x"67800000",
        2723 => x"9308d005",
        2724 => x"73000000",
        2725 => x"63520502",
        2726 => x"130101ff",
        2727 => x"23248100",
        2728 => x"13040500",
        2729 => x"23261100",
        2730 => x"33048040",
        2731 => x"efe05fc6",
        2732 => x"23208500",
        2733 => x"6f000000",
        2734 => x"6f000000",
        2735 => x"130101ff",
        2736 => x"23261100",
        2737 => x"23248100",
        2738 => x"9308900a",
        2739 => x"73000000",
        2740 => x"13040500",
        2741 => x"635a0500",
        2742 => x"33048040",
        2743 => x"efe05fc3",
        2744 => x"23208500",
        2745 => x"1304f0ff",
        2746 => x"8320c100",
        2747 => x"13050400",
        2748 => x"03248100",
        2749 => x"13010101",
        2750 => x"67800000",
        2751 => x"83a70189",
        2752 => x"130101ff",
        2753 => x"23261100",
        2754 => x"93060500",
        2755 => x"13870189",
        2756 => x"639c0702",
        2757 => x"9308600d",
        2758 => x"13050000",
        2759 => x"73000000",
        2760 => x"9307f0ff",
        2761 => x"6310f502",
        2762 => x"efe09fbe",
        2763 => x"9307c000",
        2764 => x"2320f500",
        2765 => x"1305f0ff",
        2766 => x"8320c100",
        2767 => x"13010101",
        2768 => x"67800000",
        2769 => x"2320a700",
        2770 => x"83270700",
        2771 => x"9308600d",
        2772 => x"b386f600",
        2773 => x"13850600",
        2774 => x"73000000",
        2775 => x"e316d5fc",
        2776 => x"2320a700",
        2777 => x"13850700",
        2778 => x"6ff01ffd",
        2779 => x"10000000",
        2780 => x"00000000",
        2781 => x"037a5200",
        2782 => x"017c0101",
        2783 => x"1b0d0200",
        2784 => x"10000000",
        2785 => x"18000000",
        2786 => x"c4dbffff",
        2787 => x"78040000",
        2788 => x"00000000",
        2789 => x"10000000",
        2790 => x"00000000",
        2791 => x"037a5200",
        2792 => x"017c0101",
        2793 => x"1b0d0200",
        2794 => x"10000000",
        2795 => x"18000000",
        2796 => x"14e0ffff",
        2797 => x"30040000",
        2798 => x"00000000",
        2799 => x"10000000",
        2800 => x"00000000",
        2801 => x"037a5200",
        2802 => x"017c0101",
        2803 => x"1b0d0200",
        2804 => x"10000000",
        2805 => x"18000000",
        2806 => x"1ce4ffff",
        2807 => x"e4030000",
        2808 => x"00000000",
        2809 => x"2c020000",
        2810 => x"9c010000",
        2811 => x"9c010000",
        2812 => x"9c010000",
        2813 => x"9c010000",
        2814 => x"10020000",
        2815 => x"9c010000",
        2816 => x"d0010000",
        2817 => x"9c010000",
        2818 => x"9c010000",
        2819 => x"d0010000",
        2820 => x"9c010000",
        2821 => x"9c010000",
        2822 => x"9c010000",
        2823 => x"9c010000",
        2824 => x"9c010000",
        2825 => x"9c010000",
        2826 => x"9c010000",
        2827 => x"80010000",
        2828 => x"28040000",
        2829 => x"28040000",
        2830 => x"28040000",
        2831 => x"80040000",
        2832 => x"28040000",
        2833 => x"28040000",
        2834 => x"28040000",
        2835 => x"28040000",
        2836 => x"28040000",
        2837 => x"28040000",
        2838 => x"28040000",
        2839 => x"48040000",
        2840 => x"ec040000",
        2841 => x"b4040000",
        2842 => x"b4040000",
        2843 => x"b4040000",
        2844 => x"b4040000",
        2845 => x"e0040000",
        2846 => x"74050000",
        2847 => x"4c050000",
        2848 => x"b4040000",
        2849 => x"b4040000",
        2850 => x"b4040000",
        2851 => x"b4040000",
        2852 => x"b4040000",
        2853 => x"b4040000",
        2854 => x"b4040000",
        2855 => x"b4040000",
        2856 => x"b4040000",
        2857 => x"b4040000",
        2858 => x"b4040000",
        2859 => x"b4040000",
        2860 => x"b4040000",
        2861 => x"b4040000",
        2862 => x"cc040000",
        2863 => x"cc040000",
        2864 => x"b4040000",
        2865 => x"b4040000",
        2866 => x"b4040000",
        2867 => x"b4040000",
        2868 => x"b4040000",
        2869 => x"b4040000",
        2870 => x"b4040000",
        2871 => x"b4040000",
        2872 => x"b4040000",
        2873 => x"b4040000",
        2874 => x"b4040000",
        2875 => x"b4040000",
        2876 => x"e0040000",
        2877 => x"ec040000",
        2878 => x"04050000",
        2879 => x"34050000",
        2880 => x"b4040000",
        2881 => x"b4040000",
        2882 => x"b4040000",
        2883 => x"b4040000",
        2884 => x"b4040000",
        2885 => x"b4040000",
        2886 => x"1c050000",
        2887 => x"b4040000",
        2888 => x"b4040000",
        2889 => x"b4040000",
        2890 => x"b4040000",
        2891 => x"cc040000",
        2892 => x"cc040000",
        2893 => x"00010202",
        2894 => x"03030303",
        2895 => x"04040404",
        2896 => x"04040404",
        2897 => x"05050505",
        2898 => x"05050505",
        2899 => x"05050505",
        2900 => x"05050505",
        2901 => x"06060606",
        2902 => x"06060606",
        2903 => x"06060606",
        2904 => x"06060606",
        2905 => x"06060606",
        2906 => x"06060606",
        2907 => x"06060606",
        2908 => x"06060606",
        2909 => x"07070707",
        2910 => x"07070707",
        2911 => x"07070707",
        2912 => x"07070707",
        2913 => x"07070707",
        2914 => x"07070707",
        2915 => x"07070707",
        2916 => x"07070707",
        2917 => x"07070707",
        2918 => x"07070707",
        2919 => x"07070707",
        2920 => x"07070707",
        2921 => x"07070707",
        2922 => x"07070707",
        2923 => x"07070707",
        2924 => x"07070707",
        2925 => x"08080808",
        2926 => x"08080808",
        2927 => x"08080808",
        2928 => x"08080808",
        2929 => x"08080808",
        2930 => x"08080808",
        2931 => x"08080808",
        2932 => x"08080808",
        2933 => x"08080808",
        2934 => x"08080808",
        2935 => x"08080808",
        2936 => x"08080808",
        2937 => x"08080808",
        2938 => x"08080808",
        2939 => x"08080808",
        2940 => x"08080808",
        2941 => x"08080808",
        2942 => x"08080808",
        2943 => x"08080808",
        2944 => x"08080808",
        2945 => x"08080808",
        2946 => x"08080808",
        2947 => x"08080808",
        2948 => x"08080808",
        2949 => x"08080808",
        2950 => x"08080808",
        2951 => x"08080808",
        2952 => x"08080808",
        2953 => x"08080808",
        2954 => x"08080808",
        2955 => x"08080808",
        2956 => x"08080808",
        2957 => x"0d0a0d0a",
        2958 => x"44697370",
        2959 => x"6c617969",
        2960 => x"6e672074",
        2961 => x"68652074",
        2962 => x"696d6520",
        2963 => x"70617373",
        2964 => x"65642073",
        2965 => x"696e6365",
        2966 => x"20726573",
        2967 => x"65740d0a",
        2968 => x"0d0a0000",
        2969 => x"2530356c",
        2970 => x"643a2530",
        2971 => x"366c6420",
        2972 => x"20202530",
        2973 => x"326c643a",
        2974 => x"2530326c",
        2975 => x"643a2530",
        2976 => x"326c640d",
        2977 => x"00000000",
        2978 => x"696e7465",
        2979 => x"72727570",
        2980 => x"745f6469",
        2981 => x"72656374",
        2982 => x"00000000",
        2983 => x"52495343",
        2984 => x"2d562052",
        2985 => x"56333249",
        2986 => x"4d206261",
        2987 => x"7265206d",
        2988 => x"6574616c",
        2989 => x"2070726f",
        2990 => x"63657373",
        2991 => x"6f720000",
        2992 => x"54686520",
        2993 => x"48616775",
        2994 => x"6520556e",
        2995 => x"69766572",
        2996 => x"73697479",
        2997 => x"206f6620",
        2998 => x"4170706c",
        2999 => x"69656420",
        3000 => x"53636965",
        3001 => x"6e636573",
        3002 => x"00000000",
        3003 => x"44657061",
        3004 => x"72746d65",
        3005 => x"6e74206f",
        3006 => x"6620456c",
        3007 => x"65637472",
        3008 => x"6963616c",
        3009 => x"20456e67",
        3010 => x"696e6565",
        3011 => x"72696e67",
        3012 => x"00000000",
        3013 => x"4a2e452e",
        3014 => x"4a2e206f",
        3015 => x"70206465",
        3016 => x"6e204272",
        3017 => x"6f757700",
        3018 => x"3c627265",
        3019 => x"616b3e0d",
        3020 => x"0a000000",
        3021 => x"0d0a4542",
        3022 => x"5245414b",
        3023 => x"21206d69",
        3024 => x"70203d20",
        3025 => x"00000000",
        3026 => x"232d302b",
        3027 => x"20000000",
        3028 => x"686c4c00",
        3029 => x"65666745",
        3030 => x"46470000",
        3031 => x"30313233",
        3032 => x"34353637",
        3033 => x"38394142",
        3034 => x"43444546",
        3035 => x"00000000",
        3036 => x"30313233",
        3037 => x"34353637",
        3038 => x"38396162",
        3039 => x"63646566",
        3040 => x"00000000",
        3041 => x"30220000",
        3042 => x"50220000",
        3043 => x"fc210000",
        3044 => x"fc210000",
        3045 => x"fc210000",
        3046 => x"fc210000",
        3047 => x"50220000",
        3048 => x"fc210000",
        3049 => x"fc210000",
        3050 => x"fc210000",
        3051 => x"fc210000",
        3052 => x"3c240000",
        3053 => x"a8220000",
        3054 => x"b8230000",
        3055 => x"fc210000",
        3056 => x"fc210000",
        3057 => x"84240000",
        3058 => x"fc210000",
        3059 => x"a8220000",
        3060 => x"fc210000",
        3061 => x"fc210000",
        3062 => x"c4230000",
        3063 => x"18000020",
        3064 => x"882e0000",
        3065 => x"9c2e0000",
        3066 => x"c02e0000",
        3067 => x"ec2e0000",
        3068 => x"142f0000",
        3069 => x"00000000",
        3070 => x"00000000",
        3071 => x"00000000",
        3072 => x"00000000",
        3073 => x"00000000",
        3074 => x"00000000",
        3075 => x"00000000",
        3076 => x"00000000",
        3077 => x"00000000",
        3078 => x"00000000",
        3079 => x"00000000",
        3080 => x"00000000",
        3081 => x"00000000",
        3082 => x"00000000",
        3083 => x"00000000",
        3084 => x"00000000",
        3085 => x"00000000",
        3086 => x"00000000",
        3087 => x"00000000",
        3088 => x"00000000",
        3089 => x"00000000",
        3090 => x"00000000",
        3091 => x"00000000",
        3092 => x"00000000",
        3093 => x"00000000",
        3094 => x"80000020",
        3095 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
