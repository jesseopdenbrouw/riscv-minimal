-- srec2vhdl table generator
-- for input file flash.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97",    1 => x"11",    2 => x"00",    3 => x"20", 
           4 => x"93",    5 => x"81",    6 => x"01",    7 => x"80", 
           8 => x"17",    9 => x"41",   10 => x"00",   11 => x"20", 
          12 => x"13",   13 => x"01",   14 => x"81",   15 => x"ff", 
          16 => x"97",   17 => x"00",   18 => x"00",   19 => x"00", 
          20 => x"e7",   21 => x"80",   22 => x"c0",   23 => x"00", 
          24 => x"6f",   25 => x"00",   26 => x"00",   27 => x"00", 
          28 => x"b7",   29 => x"06",   30 => x"00",   31 => x"f0", 
          32 => x"37",   33 => x"57",   34 => x"4c",   35 => x"00", 
          36 => x"13",   37 => x"01",   38 => x"01",   39 => x"ff", 
          40 => x"93",   41 => x"86",   42 => x"46",   43 => x"00", 
          44 => x"13",   45 => x"06",   46 => x"f0",   47 => x"ff", 
          48 => x"13",   49 => x"07",   50 => x"f7",   51 => x"b3", 
          52 => x"23",   53 => x"a0",   54 => x"c6",   55 => x"00", 
          56 => x"23",   57 => x"26",   58 => x"01",   59 => x"00", 
          60 => x"83",   61 => x"27",   62 => x"c1",   63 => x"00", 
          64 => x"63",   65 => x"6c",   66 => x"f7",   67 => x"00", 
          68 => x"83",   69 => x"27",   70 => x"c1",   71 => x"00", 
          72 => x"93",   73 => x"87",   74 => x"17",   75 => x"00", 
          76 => x"23",   77 => x"26",   78 => x"f1",   79 => x"00", 
          80 => x"83",   81 => x"27",   82 => x"c1",   83 => x"00", 
          84 => x"e3",   85 => x"78",   86 => x"f7",   87 => x"fe", 
          88 => x"83",   89 => x"a7",   90 => x"06",   91 => x"00", 
          92 => x"93",   93 => x"c7",   94 => x"f7",   95 => x"ff", 
          96 => x"23",   97 => x"a0",   98 => x"f6",   99 => x"00", 
         100 => x"23",  101 => x"26",  102 => x"01",  103 => x"00", 
         104 => x"83",  105 => x"27",  106 => x"c1",  107 => x"00", 
         108 => x"e3",  109 => x"64",  110 => x"f7",  111 => x"fc", 
         112 => x"83",  113 => x"27",  114 => x"c1",  115 => x"00", 
         116 => x"93",  117 => x"87",  118 => x"17",  119 => x"00", 
         120 => x"23",  121 => x"26",  122 => x"f1",  123 => x"00", 
         124 => x"83",  125 => x"27",  126 => x"c1",  127 => x"00", 
         128 => x"e3",  129 => x"78",  130 => x"f7",  131 => x"fe", 
         132 => x"6f",  133 => x"f0",  134 => x"1f",  135 => x"fb", 
        others => (others => '-')
    );
end package processor_common_rom;
