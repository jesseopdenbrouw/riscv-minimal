-- srec2vhdl table generator
-- for input file interval.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"13874186",
           5 => x"93864187",
           6 => x"637ed700",
           7 => x"93874186",
           8 => x"23800700",
           9 => x"13870700",
          10 => x"03470700",
          11 => x"93871700",
          12 => x"e398d7fe",
          13 => x"b7070020",
          14 => x"13870700",
          15 => x"13864186",
          16 => x"6374c702",
          17 => x"b7260000",
          18 => x"93860680",
          19 => x"93870700",
          20 => x"03c70600",
          21 => x"93871700",
          22 => x"93861600",
          23 => x"1377f70f",
          24 => x"a38fe7fe",
          25 => x"e396c7fe",
          26 => x"ef008033",
          27 => x"ef00001c",
          28 => x"ef008017",
          29 => x"83470500",
          30 => x"63820702",
          31 => x"370700f0",
          32 => x"13051500",
          33 => x"2320f702",
          34 => x"8327c702",
          35 => x"93f70701",
          36 => x"e38c07fe",
          37 => x"83470500",
          38 => x"e39407fe",
          39 => x"67800000",
          40 => x"37170000",
          41 => x"b70700f0",
          42 => x"13077745",
          43 => x"23a2e702",
          44 => x"67800000",
          45 => x"1375f50f",
          46 => x"b70700f0",
          47 => x"23a0a702",
          48 => x"370700f0",
          49 => x"8327c702",
          50 => x"93f70701",
          51 => x"e38c07fe",
          52 => x"67800000",
          53 => x"63060502",
          54 => x"83470500",
          55 => x"63820702",
          56 => x"370700f0",
          57 => x"13051500",
          58 => x"2320f702",
          59 => x"8327c702",
          60 => x"93f70701",
          61 => x"e38c07fe",
          62 => x"83470500",
          63 => x"e39407fe",
          64 => x"67800000",
          65 => x"13030500",
          66 => x"630a0600",
          67 => x"2300b300",
          68 => x"1306f6ff",
          69 => x"13031300",
          70 => x"e31a06fe",
          71 => x"67800000",
          72 => x"13030500",
          73 => x"630e0600",
          74 => x"83830500",
          75 => x"23007300",
          76 => x"1306f6ff",
          77 => x"13031300",
          78 => x"93851500",
          79 => x"e31606fe",
          80 => x"67800000",
          81 => x"630c0602",
          82 => x"13030500",
          83 => x"93061000",
          84 => x"636ab500",
          85 => x"9306f0ff",
          86 => x"1307f6ff",
          87 => x"3303e300",
          88 => x"b385e500",
          89 => x"83830500",
          90 => x"23007300",
          91 => x"1306f6ff",
          92 => x"3303d300",
          93 => x"b385d500",
          94 => x"e31606fe",
          95 => x"67800000",
          96 => x"03a74186",
          97 => x"b7870020",
          98 => x"93870700",
          99 => x"93060040",
         100 => x"b387d740",
         101 => x"630c0700",
         102 => x"3305a700",
         103 => x"63e2a702",
         104 => x"23a2a186",
         105 => x"13050700",
         106 => x"67800000",
         107 => x"93868187",
         108 => x"13878187",
         109 => x"23a2d186",
         110 => x"3305a700",
         111 => x"e3f2a7fe",
         112 => x"130101ff",
         113 => x"23261100",
         114 => x"ef00c005",
         115 => x"8320c100",
         116 => x"9307c000",
         117 => x"2320f500",
         118 => x"1307f0ff",
         119 => x"13050700",
         120 => x"13010101",
         121 => x"67800000",
         122 => x"6f000000",
         123 => x"93070000",
         124 => x"13070500",
         125 => x"93860700",
         126 => x"13860700",
         127 => x"f32710c8",
         128 => x"f32610c0",
         129 => x"732610c8",
         130 => x"e39ac7fe",
         131 => x"13050000",
         132 => x"2320d700",
         133 => x"23220700",
         134 => x"23240700",
         135 => x"23260700",
         136 => x"67800000",
         137 => x"03a50186",
         138 => x"67800000",
         139 => x"130101f7",
         140 => x"13060006",
         141 => x"93050000",
         142 => x"13050101",
         143 => x"23261108",
         144 => x"23248108",
         145 => x"23229108",
         146 => x"23202109",
         147 => x"232e3107",
         148 => x"232c4107",
         149 => x"232a5107",
         150 => x"23260100",
         151 => x"eff09fea",
         152 => x"37170000",
         153 => x"b70700f0",
         154 => x"13077745",
         155 => x"37150000",
         156 => x"23a2e702",
         157 => x"13050573",
         158 => x"eff0dfdf",
         159 => x"b7460f00",
         160 => x"37160000",
         161 => x"93860624",
         162 => x"13068674",
         163 => x"93054006",
         164 => x"1305c100",
         165 => x"ef00c025",
         166 => x"1305c100",
         167 => x"b7190000",
         168 => x"37190000",
         169 => x"b7544c00",
         170 => x"eff0dfdc",
         171 => x"371a0000",
         172 => x"93890971",
         173 => x"1309c971",
         174 => x"370400f0",
         175 => x"9384f4b3",
         176 => x"ef00c009",
         177 => x"93060500",
         178 => x"930a0500",
         179 => x"13060a76",
         180 => x"93054006",
         181 => x"1305c100",
         182 => x"ef008021",
         183 => x"8347c100",
         184 => x"63820702",
         185 => x"1307c100",
         186 => x"13071700",
         187 => x"2320f402",
         188 => x"8327c402",
         189 => x"93f70701",
         190 => x"e38c07fe",
         191 => x"83470700",
         192 => x"e39407fe",
         193 => x"93077005",
         194 => x"13870900",
         195 => x"13071700",
         196 => x"2320f402",
         197 => x"8327c402",
         198 => x"93f70701",
         199 => x"e38c07fe",
         200 => x"83470700",
         201 => x"e39407fe",
         202 => x"ef004003",
         203 => x"33055541",
         204 => x"e3fca4fe",
         205 => x"93075003",
         206 => x"13070900",
         207 => x"13071700",
         208 => x"2320f402",
         209 => x"8327c402",
         210 => x"93f70701",
         211 => x"e38c07fe",
         212 => x"83470700",
         213 => x"e39407fe",
         214 => x"6ff09ff6",
         215 => x"03a50186",
         216 => x"130101fe",
         217 => x"93050100",
         218 => x"232e1100",
         219 => x"ef008023",
         220 => x"9307f0ff",
         221 => x"6300f502",
         222 => x"83274100",
         223 => x"03250100",
         224 => x"3305f500",
         225 => x"83278100",
         226 => x"3305f500",
         227 => x"8327c100",
         228 => x"3305f500",
         229 => x"8320c101",
         230 => x"13010102",
         231 => x"67800000",
         232 => x"130101ff",
         233 => x"23248100",
         234 => x"23229100",
         235 => x"37240000",
         236 => x"b7240000",
         237 => x"93870480",
         238 => x"13040480",
         239 => x"3304f440",
         240 => x"23202101",
         241 => x"23261100",
         242 => x"13542440",
         243 => x"93840480",
         244 => x"13090000",
         245 => x"63108904",
         246 => x"b7240000",
         247 => x"37240000",
         248 => x"93870480",
         249 => x"13040480",
         250 => x"3304f440",
         251 => x"13542440",
         252 => x"93840480",
         253 => x"13090000",
         254 => x"63188902",
         255 => x"8320c100",
         256 => x"03248100",
         257 => x"83244100",
         258 => x"03290100",
         259 => x"13010101",
         260 => x"67800000",
         261 => x"83a70400",
         262 => x"13091900",
         263 => x"93844400",
         264 => x"e7800700",
         265 => x"6ff01ffb",
         266 => x"83a70400",
         267 => x"13091900",
         268 => x"93844400",
         269 => x"e7800700",
         270 => x"6ff01ffc",
         271 => x"130101f7",
         272 => x"232c8106",
         273 => x"232a9106",
         274 => x"232e1106",
         275 => x"23282107",
         276 => x"2320e108",
         277 => x"2322f108",
         278 => x"23240109",
         279 => x"23261109",
         280 => x"93040500",
         281 => x"13040600",
         282 => x"63540602",
         283 => x"9307b008",
         284 => x"2320f500",
         285 => x"1305f0ff",
         286 => x"8320c107",
         287 => x"03248107",
         288 => x"83244107",
         289 => x"03290107",
         290 => x"13010109",
         291 => x"67800000",
         292 => x"93078020",
         293 => x"231af100",
         294 => x"2324b100",
         295 => x"232cb100",
         296 => x"13860600",
         297 => x"93070000",
         298 => x"63040400",
         299 => x"9307f4ff",
         300 => x"1309f0ff",
         301 => x"93060108",
         302 => x"93058100",
         303 => x"13850400",
         304 => x"2328f100",
         305 => x"232ef100",
         306 => x"231b2101",
         307 => x"2322d100",
         308 => x"ef00c040",
         309 => x"63562501",
         310 => x"9307b008",
         311 => x"23a0f400",
         312 => x"e30c04f8",
         313 => x"83278100",
         314 => x"23800700",
         315 => x"6ff0dff8",
         316 => x"130101f6",
         317 => x"232a9106",
         318 => x"232af108",
         319 => x"232e1106",
         320 => x"232c8106",
         321 => x"23282107",
         322 => x"2326d108",
         323 => x"2328e108",
         324 => x"232c0109",
         325 => x"232e1109",
         326 => x"83a40186",
         327 => x"63d40502",
         328 => x"9307b008",
         329 => x"23a0f400",
         330 => x"1305f0ff",
         331 => x"8320c107",
         332 => x"03248107",
         333 => x"83244107",
         334 => x"03290107",
         335 => x"1301010a",
         336 => x"67800000",
         337 => x"93078020",
         338 => x"231af100",
         339 => x"2324a100",
         340 => x"232ca100",
         341 => x"13840500",
         342 => x"93070000",
         343 => x"63840500",
         344 => x"9387f5ff",
         345 => x"1309f0ff",
         346 => x"9306c108",
         347 => x"93058100",
         348 => x"13850400",
         349 => x"2328f100",
         350 => x"232ef100",
         351 => x"231b2101",
         352 => x"2322d100",
         353 => x"ef008035",
         354 => x"63562501",
         355 => x"9307b008",
         356 => x"23a0f400",
         357 => x"e30c04f8",
         358 => x"83278100",
         359 => x"23800700",
         360 => x"6ff0dff8",
         361 => x"13850500",
         362 => x"6ff05fc4",
         363 => x"130101fe",
         364 => x"23282101",
         365 => x"03a98500",
         366 => x"232c8100",
         367 => x"23263101",
         368 => x"23244101",
         369 => x"23225101",
         370 => x"232e1100",
         371 => x"232a9100",
         372 => x"23206101",
         373 => x"83aa0500",
         374 => x"13840500",
         375 => x"130a0600",
         376 => x"93890600",
         377 => x"63ec2609",
         378 => x"83d7c500",
         379 => x"13f70748",
         380 => x"63040708",
         381 => x"03274401",
         382 => x"93043000",
         383 => x"83a50501",
         384 => x"b384e402",
         385 => x"13072000",
         386 => x"b38aba40",
         387 => x"130b0500",
         388 => x"b3c4e402",
         389 => x"13871600",
         390 => x"33075701",
         391 => x"63f4e400",
         392 => x"93040700",
         393 => x"93f70740",
         394 => x"6386070a",
         395 => x"93850400",
         396 => x"13050b00",
         397 => x"ef00504a",
         398 => x"13090500",
         399 => x"630c050a",
         400 => x"83250401",
         401 => x"13860a00",
         402 => x"eff09fad",
         403 => x"8357c400",
         404 => x"93f7f7b7",
         405 => x"93e70708",
         406 => x"2316f400",
         407 => x"23282401",
         408 => x"232a9400",
         409 => x"33095901",
         410 => x"b3845441",
         411 => x"23202401",
         412 => x"23249400",
         413 => x"13890900",
         414 => x"63f42901",
         415 => x"13890900",
         416 => x"03250400",
         417 => x"13060900",
         418 => x"93050a00",
         419 => x"eff09fab",
         420 => x"83278400",
         421 => x"13050000",
         422 => x"b3872741",
         423 => x"2324f400",
         424 => x"83270400",
         425 => x"b3872701",
         426 => x"2320f400",
         427 => x"8320c101",
         428 => x"03248101",
         429 => x"83244101",
         430 => x"03290101",
         431 => x"8329c100",
         432 => x"032a8100",
         433 => x"832a4100",
         434 => x"032b0100",
         435 => x"13010102",
         436 => x"67800000",
         437 => x"13860400",
         438 => x"13050b00",
         439 => x"ef00d054",
         440 => x"13090500",
         441 => x"e31c05f6",
         442 => x"83250401",
         443 => x"13050b00",
         444 => x"ef00102f",
         445 => x"9307c000",
         446 => x"2320fb00",
         447 => x"8357c400",
         448 => x"1305f0ff",
         449 => x"93e70704",
         450 => x"2316f400",
         451 => x"6ff01ffa",
         452 => x"83278600",
         453 => x"130101fd",
         454 => x"232e3101",
         455 => x"23286101",
         456 => x"23261102",
         457 => x"23248102",
         458 => x"23229102",
         459 => x"23202103",
         460 => x"232c4101",
         461 => x"232a5101",
         462 => x"23267101",
         463 => x"23248101",
         464 => x"23229101",
         465 => x"2320a101",
         466 => x"032b0600",
         467 => x"93090600",
         468 => x"63980712",
         469 => x"13050000",
         470 => x"8320c102",
         471 => x"03248102",
         472 => x"23a20900",
         473 => x"83244102",
         474 => x"03290102",
         475 => x"8329c101",
         476 => x"032a8101",
         477 => x"832a4101",
         478 => x"032b0101",
         479 => x"832bc100",
         480 => x"032c8100",
         481 => x"832c4100",
         482 => x"032d0100",
         483 => x"13010103",
         484 => x"67800000",
         485 => x"832a0b00",
         486 => x"032d4b00",
         487 => x"130b8b00",
         488 => x"03298400",
         489 => x"832c0400",
         490 => x"e3060dfe",
         491 => x"63642d09",
         492 => x"8357c400",
         493 => x"13f70748",
         494 => x"630e0706",
         495 => x"83244401",
         496 => x"83250401",
         497 => x"b3849b02",
         498 => x"b38cbc40",
         499 => x"13871c00",
         500 => x"3307a701",
         501 => x"b3c48403",
         502 => x"63f4e400",
         503 => x"93040700",
         504 => x"93f70740",
         505 => x"638c070a",
         506 => x"93850400",
         507 => x"13050a00",
         508 => x"ef00902e",
         509 => x"13090500",
         510 => x"6302050c",
         511 => x"83250401",
         512 => x"13860c00",
         513 => x"eff0df91",
         514 => x"8357c400",
         515 => x"93f7f7b7",
         516 => x"93e70708",
         517 => x"2316f400",
         518 => x"23282401",
         519 => x"232a9400",
         520 => x"33099901",
         521 => x"b3849441",
         522 => x"23202401",
         523 => x"23249400",
         524 => x"13090d00",
         525 => x"63742d01",
         526 => x"13090d00",
         527 => x"03250400",
         528 => x"93850a00",
         529 => x"13060900",
         530 => x"eff0df8f",
         531 => x"83278400",
         532 => x"b38aaa01",
         533 => x"b3872741",
         534 => x"2324f400",
         535 => x"83270400",
         536 => x"b3872701",
         537 => x"2320f400",
         538 => x"83a78900",
         539 => x"b387a741",
         540 => x"23a4f900",
         541 => x"e38007ee",
         542 => x"130d0000",
         543 => x"6ff05ff2",
         544 => x"130a0500",
         545 => x"13840500",
         546 => x"930a0000",
         547 => x"130d0000",
         548 => x"930b3000",
         549 => x"130c2000",
         550 => x"6ff09ff0",
         551 => x"13860400",
         552 => x"13050a00",
         553 => x"ef005038",
         554 => x"13090500",
         555 => x"e31605f6",
         556 => x"83250401",
         557 => x"13050a00",
         558 => x"ef009012",
         559 => x"9307c000",
         560 => x"2320fa00",
         561 => x"8357c400",
         562 => x"1305f0ff",
         563 => x"93e70704",
         564 => x"2316f400",
         565 => x"23a40900",
         566 => x"6ff01fe8",
         567 => x"83d7c500",
         568 => x"130101f5",
         569 => x"2324810a",
         570 => x"2322910a",
         571 => x"2320210b",
         572 => x"232c4109",
         573 => x"2326110a",
         574 => x"232e3109",
         575 => x"232a5109",
         576 => x"23286109",
         577 => x"23267109",
         578 => x"23248109",
         579 => x"23229109",
         580 => x"2320a109",
         581 => x"232eb107",
         582 => x"93f70708",
         583 => x"130a0500",
         584 => x"13890500",
         585 => x"93040600",
         586 => x"13840600",
         587 => x"63880706",
         588 => x"83a70501",
         589 => x"63940706",
         590 => x"93050004",
         591 => x"ef00d019",
         592 => x"2320a900",
         593 => x"2328a900",
         594 => x"63160504",
         595 => x"9307c000",
         596 => x"2320fa00",
         597 => x"1305f0ff",
         598 => x"8320c10a",
         599 => x"0324810a",
         600 => x"8324410a",
         601 => x"0329010a",
         602 => x"8329c109",
         603 => x"032a8109",
         604 => x"832a4109",
         605 => x"032b0109",
         606 => x"832bc108",
         607 => x"032c8108",
         608 => x"832c4108",
         609 => x"032d0108",
         610 => x"832dc107",
         611 => x"1301010b",
         612 => x"67800000",
         613 => x"93070004",
         614 => x"232af900",
         615 => x"93070002",
         616 => x"a304f102",
         617 => x"93070003",
         618 => x"23220102",
         619 => x"2305f102",
         620 => x"23268100",
         621 => x"930c5002",
         622 => x"371b0000",
         623 => x"b71b0000",
         624 => x"371d0000",
         625 => x"930a0000",
         626 => x"13840400",
         627 => x"83470400",
         628 => x"63840700",
         629 => x"639c970d",
         630 => x"b30d9440",
         631 => x"63069402",
         632 => x"93860d00",
         633 => x"13860400",
         634 => x"93050900",
         635 => x"13050a00",
         636 => x"eff0dfbb",
         637 => x"9307f0ff",
         638 => x"6306f524",
         639 => x"83274102",
         640 => x"b387b701",
         641 => x"2322f102",
         642 => x"83470400",
         643 => x"638c0722",
         644 => x"9307f0ff",
         645 => x"93041400",
         646 => x"23280100",
         647 => x"232e0100",
         648 => x"232af100",
         649 => x"232c0100",
         650 => x"a3090104",
         651 => x"23240106",
         652 => x"930d1000",
         653 => x"83c50400",
         654 => x"13065000",
         655 => x"13058b76",
         656 => x"ef00c077",
         657 => x"83270101",
         658 => x"13841400",
         659 => x"63140506",
         660 => x"13f70701",
         661 => x"63060700",
         662 => x"13070002",
         663 => x"a309e104",
         664 => x"13f78700",
         665 => x"63060700",
         666 => x"1307b002",
         667 => x"a309e104",
         668 => x"83c60400",
         669 => x"1307a002",
         670 => x"638ce604",
         671 => x"8327c101",
         672 => x"13840400",
         673 => x"93060000",
         674 => x"13069000",
         675 => x"1305a000",
         676 => x"03470400",
         677 => x"93051400",
         678 => x"130707fd",
         679 => x"637ce608",
         680 => x"63840604",
         681 => x"232ef100",
         682 => x"6f000004",
         683 => x"13041400",
         684 => x"6ff0dff1",
         685 => x"13078b76",
         686 => x"3305e540",
         687 => x"3395ad00",
         688 => x"b3e7a700",
         689 => x"2328f100",
         690 => x"93040400",
         691 => x"6ff09ff6",
         692 => x"0327c100",
         693 => x"93064700",
         694 => x"03270700",
         695 => x"2326d100",
         696 => x"63400704",
         697 => x"232ee100",
         698 => x"03470400",
         699 => x"9307e002",
         700 => x"6316f708",
         701 => x"03471400",
         702 => x"9307a002",
         703 => x"631af704",
         704 => x"8327c100",
         705 => x"13042400",
         706 => x"13874700",
         707 => x"83a70700",
         708 => x"2326e100",
         709 => x"63ca0702",
         710 => x"232af100",
         711 => x"6f000006",
         712 => x"3307e040",
         713 => x"93e72700",
         714 => x"232ee100",
         715 => x"2328f100",
         716 => x"6ff09ffb",
         717 => x"b387a702",
         718 => x"13840500",
         719 => x"93061000",
         720 => x"b387e700",
         721 => x"6ff0dff4",
         722 => x"9307f0ff",
         723 => x"6ff0dffc",
         724 => x"13041400",
         725 => x"232a0100",
         726 => x"93060000",
         727 => x"93070000",
         728 => x"13069000",
         729 => x"1305a000",
         730 => x"03470400",
         731 => x"93051400",
         732 => x"130707fd",
         733 => x"6372e608",
         734 => x"e39006fa",
         735 => x"83450400",
         736 => x"13063000",
         737 => x"13850b77",
         738 => x"ef004063",
         739 => x"63020502",
         740 => x"93870b77",
         741 => x"3305f540",
         742 => x"83270101",
         743 => x"13070004",
         744 => x"3317a700",
         745 => x"b3e7e700",
         746 => x"13041400",
         747 => x"2328f100",
         748 => x"83450400",
         749 => x"13066000",
         750 => x"13054d77",
         751 => x"93041400",
         752 => x"2304b102",
         753 => x"ef00805f",
         754 => x"630a0508",
         755 => x"63980a04",
         756 => x"03270101",
         757 => x"8327c100",
         758 => x"13770710",
         759 => x"63080702",
         760 => x"93874700",
         761 => x"2326f100",
         762 => x"83274102",
         763 => x"b3873701",
         764 => x"2322f102",
         765 => x"6ff05fdd",
         766 => x"b387a702",
         767 => x"13840500",
         768 => x"93061000",
         769 => x"b387e700",
         770 => x"6ff01ff6",
         771 => x"93877700",
         772 => x"93f787ff",
         773 => x"93878700",
         774 => x"6ff0dffc",
         775 => x"1307c100",
         776 => x"9306c05a",
         777 => x"13060900",
         778 => x"93050101",
         779 => x"13050a00",
         780 => x"97000000",
         781 => x"e7000000",
         782 => x"9307f0ff",
         783 => x"93090500",
         784 => x"e314f5fa",
         785 => x"8357c900",
         786 => x"1305f0ff",
         787 => x"93f70704",
         788 => x"e39407d0",
         789 => x"03254102",
         790 => x"6ff01fd0",
         791 => x"1307c100",
         792 => x"9306c05a",
         793 => x"13060900",
         794 => x"93050101",
         795 => x"13050a00",
         796 => x"ef00801b",
         797 => x"6ff05ffc",
         798 => x"130101fd",
         799 => x"232c4101",
         800 => x"83a70501",
         801 => x"130a0700",
         802 => x"03a78500",
         803 => x"23248102",
         804 => x"23202103",
         805 => x"232e3101",
         806 => x"232a5101",
         807 => x"23261102",
         808 => x"23229102",
         809 => x"23286101",
         810 => x"23267101",
         811 => x"93090500",
         812 => x"13840500",
         813 => x"13090600",
         814 => x"938a0600",
         815 => x"63d4e700",
         816 => x"93070700",
         817 => x"2320f900",
         818 => x"03473404",
         819 => x"63060700",
         820 => x"93871700",
         821 => x"2320f900",
         822 => x"83270400",
         823 => x"93f70702",
         824 => x"63880700",
         825 => x"83270900",
         826 => x"93872700",
         827 => x"2320f900",
         828 => x"83240400",
         829 => x"93f46400",
         830 => x"639e0400",
         831 => x"130b9401",
         832 => x"930bf0ff",
         833 => x"8327c400",
         834 => x"03270900",
         835 => x"b387e740",
         836 => x"63c2f408",
         837 => x"83473404",
         838 => x"b336f000",
         839 => x"83270400",
         840 => x"93f70702",
         841 => x"6390070c",
         842 => x"13063404",
         843 => x"93850a00",
         844 => x"13850900",
         845 => x"e7000a00",
         846 => x"9307f0ff",
         847 => x"6308f506",
         848 => x"83270400",
         849 => x"13074000",
         850 => x"93040000",
         851 => x"93f76700",
         852 => x"639ce700",
         853 => x"8324c400",
         854 => x"83270900",
         855 => x"b384f440",
         856 => x"63d40400",
         857 => x"93040000",
         858 => x"83278400",
         859 => x"03270401",
         860 => x"6356f700",
         861 => x"b387e740",
         862 => x"b384f400",
         863 => x"13090000",
         864 => x"1304a401",
         865 => x"130bf0ff",
         866 => x"63902409",
         867 => x"13050000",
         868 => x"6f000002",
         869 => x"93061000",
         870 => x"13060b00",
         871 => x"93850a00",
         872 => x"13850900",
         873 => x"e7000a00",
         874 => x"631a7503",
         875 => x"1305f0ff",
         876 => x"8320c102",
         877 => x"03248102",
         878 => x"83244102",
         879 => x"03290102",
         880 => x"8329c101",
         881 => x"032a8101",
         882 => x"832a4101",
         883 => x"032b0101",
         884 => x"832bc100",
         885 => x"13010103",
         886 => x"67800000",
         887 => x"93841400",
         888 => x"6ff05ff2",
         889 => x"3307d400",
         890 => x"13060003",
         891 => x"a301c704",
         892 => x"03475404",
         893 => x"93871600",
         894 => x"b307f400",
         895 => x"93862600",
         896 => x"a381e704",
         897 => x"6ff05ff2",
         898 => x"93061000",
         899 => x"13060400",
         900 => x"93850a00",
         901 => x"13850900",
         902 => x"e7000a00",
         903 => x"e30865f9",
         904 => x"13091900",
         905 => x"6ff05ff6",
         906 => x"130101fd",
         907 => x"23248102",
         908 => x"23229102",
         909 => x"23202103",
         910 => x"232e3101",
         911 => x"23261102",
         912 => x"232c4101",
         913 => x"232a5101",
         914 => x"23286101",
         915 => x"83c88501",
         916 => x"93078007",
         917 => x"93040500",
         918 => x"13840500",
         919 => x"13090600",
         920 => x"93890600",
         921 => x"63ee1701",
         922 => x"93072006",
         923 => x"93863504",
         924 => x"63ee1701",
         925 => x"63840828",
         926 => x"93078005",
         927 => x"6388f822",
         928 => x"930a2404",
         929 => x"23011405",
         930 => x"6f004004",
         931 => x"9387d8f9",
         932 => x"93f7f70f",
         933 => x"13065001",
         934 => x"e364f6fe",
         935 => x"37160000",
         936 => x"93972700",
         937 => x"1306467a",
         938 => x"b387c700",
         939 => x"83a70700",
         940 => x"67800700",
         941 => x"83270700",
         942 => x"938a2504",
         943 => x"93864700",
         944 => x"83a70700",
         945 => x"2320d700",
         946 => x"2381f504",
         947 => x"93071000",
         948 => x"6f008026",
         949 => x"83a70500",
         950 => x"03250700",
         951 => x"13f60708",
         952 => x"93054500",
         953 => x"63060602",
         954 => x"83270500",
         955 => x"2320b700",
         956 => x"37180000",
         957 => x"63d80700",
         958 => x"1307d002",
         959 => x"b307f040",
         960 => x"a301e404",
         961 => x"1308c877",
         962 => x"1307a000",
         963 => x"6f008006",
         964 => x"13f60704",
         965 => x"83270500",
         966 => x"2320b700",
         967 => x"e30a06fc",
         968 => x"93970701",
         969 => x"93d70741",
         970 => x"6ff09ffc",
         971 => x"03a60500",
         972 => x"83270700",
         973 => x"13750608",
         974 => x"93854700",
         975 => x"63080500",
         976 => x"2320b700",
         977 => x"83a70700",
         978 => x"6f004001",
         979 => x"13760604",
         980 => x"2320b700",
         981 => x"e30806fe",
         982 => x"83d70700",
         983 => x"37180000",
         984 => x"1307f006",
         985 => x"1308c877",
         986 => x"6388e814",
         987 => x"1307a000",
         988 => x"a3010404",
         989 => x"03264400",
         990 => x"2324c400",
         991 => x"63480600",
         992 => x"83250400",
         993 => x"93f5b5ff",
         994 => x"2320b400",
         995 => x"63960700",
         996 => x"938a0600",
         997 => x"63040602",
         998 => x"938a0600",
         999 => x"33f6e702",
        1000 => x"938afaff",
        1001 => x"3306c800",
        1002 => x"03460600",
        1003 => x"2380ca00",
        1004 => x"13860700",
        1005 => x"b3d7e702",
        1006 => x"e372e6fe",
        1007 => x"93078000",
        1008 => x"6314f702",
        1009 => x"83270400",
        1010 => x"93f71700",
        1011 => x"638e0700",
        1012 => x"03274400",
        1013 => x"83270401",
        1014 => x"63c8e700",
        1015 => x"93070003",
        1016 => x"a38ffafe",
        1017 => x"938afaff",
        1018 => x"b3865641",
        1019 => x"2328d400",
        1020 => x"13870900",
        1021 => x"93060900",
        1022 => x"1306c100",
        1023 => x"93050400",
        1024 => x"13850400",
        1025 => x"eff05fc7",
        1026 => x"130af0ff",
        1027 => x"631c4513",
        1028 => x"1305f0ff",
        1029 => x"8320c102",
        1030 => x"03248102",
        1031 => x"83244102",
        1032 => x"03290102",
        1033 => x"8329c101",
        1034 => x"032a8101",
        1035 => x"832a4101",
        1036 => x"032b0101",
        1037 => x"13010103",
        1038 => x"67800000",
        1039 => x"83a70500",
        1040 => x"93e70702",
        1041 => x"23a0f500",
        1042 => x"37180000",
        1043 => x"93088007",
        1044 => x"13080879",
        1045 => x"a3021405",
        1046 => x"03260400",
        1047 => x"83250700",
        1048 => x"13750608",
        1049 => x"83a70500",
        1050 => x"93854500",
        1051 => x"631a0500",
        1052 => x"13750604",
        1053 => x"63060500",
        1054 => x"93970701",
        1055 => x"93d70701",
        1056 => x"2320b700",
        1057 => x"13771600",
        1058 => x"63060700",
        1059 => x"13660602",
        1060 => x"2320c400",
        1061 => x"13070001",
        1062 => x"e39c07ec",
        1063 => x"03260400",
        1064 => x"1376f6fd",
        1065 => x"2320c400",
        1066 => x"6ff09fec",
        1067 => x"37180000",
        1068 => x"1308c877",
        1069 => x"6ff01ffa",
        1070 => x"13078000",
        1071 => x"6ff05feb",
        1072 => x"03a60500",
        1073 => x"83270700",
        1074 => x"83a54501",
        1075 => x"13780608",
        1076 => x"13854700",
        1077 => x"630a0800",
        1078 => x"2320a700",
        1079 => x"83a70700",
        1080 => x"23a0b700",
        1081 => x"6f008001",
        1082 => x"2320a700",
        1083 => x"13760604",
        1084 => x"83a70700",
        1085 => x"e30606fe",
        1086 => x"2390b700",
        1087 => x"23280400",
        1088 => x"938a0600",
        1089 => x"6ff0dfee",
        1090 => x"83270700",
        1091 => x"03a64500",
        1092 => x"93050000",
        1093 => x"93864700",
        1094 => x"2320d700",
        1095 => x"83aa0700",
        1096 => x"13850a00",
        1097 => x"ef008009",
        1098 => x"63060500",
        1099 => x"33055541",
        1100 => x"2322a400",
        1101 => x"83274400",
        1102 => x"2328f400",
        1103 => x"a3010404",
        1104 => x"6ff01feb",
        1105 => x"83260401",
        1106 => x"13860a00",
        1107 => x"93050900",
        1108 => x"13850400",
        1109 => x"e7800900",
        1110 => x"e30c45eb",
        1111 => x"83270400",
        1112 => x"93f72700",
        1113 => x"63940704",
        1114 => x"8327c100",
        1115 => x"0325c400",
        1116 => x"e352f5ea",
        1117 => x"13850700",
        1118 => x"6ff0dfe9",
        1119 => x"93061000",
        1120 => x"13860a00",
        1121 => x"93050900",
        1122 => x"13850400",
        1123 => x"e7800900",
        1124 => x"e30065e9",
        1125 => x"130a1a00",
        1126 => x"8327c400",
        1127 => x"0327c100",
        1128 => x"b387e740",
        1129 => x"e34cfafc",
        1130 => x"6ff01ffc",
        1131 => x"130a0000",
        1132 => x"930a9401",
        1133 => x"130bf0ff",
        1134 => x"6ff01ffe",
        1135 => x"93f5f50f",
        1136 => x"3306c500",
        1137 => x"6316c500",
        1138 => x"13050000",
        1139 => x"67800000",
        1140 => x"83470500",
        1141 => x"e38cb7fe",
        1142 => x"13051500",
        1143 => x"6ff09ffe",
        1144 => x"638a050e",
        1145 => x"83a7c5ff",
        1146 => x"130101fe",
        1147 => x"232c8100",
        1148 => x"232e1100",
        1149 => x"1384c5ff",
        1150 => x"63d40700",
        1151 => x"3304f400",
        1152 => x"2326a100",
        1153 => x"ef000034",
        1154 => x"83a78186",
        1155 => x"0325c100",
        1156 => x"639e0700",
        1157 => x"23220400",
        1158 => x"23a48186",
        1159 => x"03248101",
        1160 => x"8320c101",
        1161 => x"13010102",
        1162 => x"6f000032",
        1163 => x"6374f402",
        1164 => x"03260400",
        1165 => x"b306c400",
        1166 => x"639ad700",
        1167 => x"83a60700",
        1168 => x"83a74700",
        1169 => x"b386c600",
        1170 => x"2320d400",
        1171 => x"2322f400",
        1172 => x"6ff09ffc",
        1173 => x"13870700",
        1174 => x"83a74700",
        1175 => x"63840700",
        1176 => x"e37af4fe",
        1177 => x"83260700",
        1178 => x"3306d700",
        1179 => x"63188602",
        1180 => x"03260400",
        1181 => x"b386c600",
        1182 => x"2320d700",
        1183 => x"3306d700",
        1184 => x"e39ec7f8",
        1185 => x"03a60700",
        1186 => x"83a74700",
        1187 => x"b306d600",
        1188 => x"2320d700",
        1189 => x"2322f700",
        1190 => x"6ff05ff8",
        1191 => x"6378c400",
        1192 => x"9307c000",
        1193 => x"2320f500",
        1194 => x"6ff05ff7",
        1195 => x"03260400",
        1196 => x"b306c400",
        1197 => x"639ad700",
        1198 => x"83a60700",
        1199 => x"83a74700",
        1200 => x"b386c600",
        1201 => x"2320d400",
        1202 => x"2322f400",
        1203 => x"23228700",
        1204 => x"6ff0dff4",
        1205 => x"67800000",
        1206 => x"130101fe",
        1207 => x"232a9100",
        1208 => x"93843500",
        1209 => x"93f4c4ff",
        1210 => x"23282101",
        1211 => x"232e1100",
        1212 => x"232c8100",
        1213 => x"23263101",
        1214 => x"93848400",
        1215 => x"9307c000",
        1216 => x"13090500",
        1217 => x"63f4f406",
        1218 => x"9304c000",
        1219 => x"63e2b406",
        1220 => x"13050900",
        1221 => x"ef000023",
        1222 => x"03a78186",
        1223 => x"93868186",
        1224 => x"13040700",
        1225 => x"631a0406",
        1226 => x"1384c186",
        1227 => x"83270400",
        1228 => x"639a0700",
        1229 => x"93050000",
        1230 => x"13050900",
        1231 => x"ef00001c",
        1232 => x"2320a400",
        1233 => x"93850400",
        1234 => x"13050900",
        1235 => x"ef00001b",
        1236 => x"9309f0ff",
        1237 => x"631a350b",
        1238 => x"9307c000",
        1239 => x"2320f900",
        1240 => x"13050900",
        1241 => x"ef00401e",
        1242 => x"6f000001",
        1243 => x"e3d004fa",
        1244 => x"9307c000",
        1245 => x"2320f900",
        1246 => x"13050000",
        1247 => x"8320c101",
        1248 => x"03248101",
        1249 => x"83244101",
        1250 => x"03290101",
        1251 => x"8329c100",
        1252 => x"13010102",
        1253 => x"67800000",
        1254 => x"83270400",
        1255 => x"b3879740",
        1256 => x"63ce0704",
        1257 => x"1306b000",
        1258 => x"637af600",
        1259 => x"2320f400",
        1260 => x"3304f400",
        1261 => x"23209400",
        1262 => x"6f000001",
        1263 => x"83274400",
        1264 => x"631a8702",
        1265 => x"23a0f600",
        1266 => x"13050900",
        1267 => x"ef00c017",
        1268 => x"1305b400",
        1269 => x"93074400",
        1270 => x"137585ff",
        1271 => x"3307f540",
        1272 => x"e30ef5f8",
        1273 => x"3304e400",
        1274 => x"b387a740",
        1275 => x"2320f400",
        1276 => x"6ff0dff8",
        1277 => x"2322f700",
        1278 => x"6ff01ffd",
        1279 => x"13070400",
        1280 => x"03244400",
        1281 => x"6ff01ff2",
        1282 => x"13043500",
        1283 => x"1374c4ff",
        1284 => x"e30285fa",
        1285 => x"b305a440",
        1286 => x"13050900",
        1287 => x"ef00000e",
        1288 => x"e31a35f9",
        1289 => x"6ff05ff3",
        1290 => x"130101fe",
        1291 => x"232c8100",
        1292 => x"232e1100",
        1293 => x"232a9100",
        1294 => x"23282101",
        1295 => x"23263101",
        1296 => x"23244101",
        1297 => x"13040600",
        1298 => x"63940502",
        1299 => x"03248101",
        1300 => x"8320c101",
        1301 => x"83244101",
        1302 => x"03290101",
        1303 => x"8329c100",
        1304 => x"032a8100",
        1305 => x"93050600",
        1306 => x"13010102",
        1307 => x"6ff0dfe6",
        1308 => x"63180602",
        1309 => x"eff0dfd6",
        1310 => x"93040000",
        1311 => x"8320c101",
        1312 => x"03248101",
        1313 => x"03290101",
        1314 => x"8329c100",
        1315 => x"032a8100",
        1316 => x"13850400",
        1317 => x"83244101",
        1318 => x"13010102",
        1319 => x"67800000",
        1320 => x"130a0500",
        1321 => x"13890500",
        1322 => x"ef00400a",
        1323 => x"93090500",
        1324 => x"63688500",
        1325 => x"93571500",
        1326 => x"93040900",
        1327 => x"e3e087fc",
        1328 => x"93050400",
        1329 => x"13050a00",
        1330 => x"eff01fe1",
        1331 => x"93040500",
        1332 => x"e30605fa",
        1333 => x"13060400",
        1334 => x"63f48900",
        1335 => x"13860900",
        1336 => x"93050900",
        1337 => x"13850400",
        1338 => x"efe09fc3",
        1339 => x"93050900",
        1340 => x"13050a00",
        1341 => x"eff0dfce",
        1342 => x"6ff05ff8",
        1343 => x"130101ff",
        1344 => x"23248100",
        1345 => x"23229100",
        1346 => x"13040500",
        1347 => x"13850500",
        1348 => x"23261100",
        1349 => x"23a80186",
        1350 => x"efe09fc6",
        1351 => x"9307f0ff",
        1352 => x"6318f500",
        1353 => x"83a70187",
        1354 => x"63840700",
        1355 => x"2320f400",
        1356 => x"8320c100",
        1357 => x"03248100",
        1358 => x"83244100",
        1359 => x"13010101",
        1360 => x"67800000",
        1361 => x"67800000",
        1362 => x"67800000",
        1363 => x"83a7c5ff",
        1364 => x"1385c7ff",
        1365 => x"63d80700",
        1366 => x"b385a500",
        1367 => x"83a70500",
        1368 => x"3305f500",
        1369 => x"67800000",
        1370 => x"130101ff",
        1371 => x"23248100",
        1372 => x"13840500",
        1373 => x"83a50500",
        1374 => x"23229100",
        1375 => x"23261100",
        1376 => x"93040500",
        1377 => x"63840500",
        1378 => x"eff01ffe",
        1379 => x"93050400",
        1380 => x"03248100",
        1381 => x"8320c100",
        1382 => x"13850400",
        1383 => x"83244100",
        1384 => x"13010101",
        1385 => x"6ff0dfc3",
        1386 => x"83a70186",
        1387 => x"6380a716",
        1388 => x"83274502",
        1389 => x"130101fe",
        1390 => x"232c8100",
        1391 => x"232e1100",
        1392 => x"232a9100",
        1393 => x"23282101",
        1394 => x"23263101",
        1395 => x"13040500",
        1396 => x"63840702",
        1397 => x"83a7c700",
        1398 => x"93040000",
        1399 => x"13090008",
        1400 => x"6392070e",
        1401 => x"83274402",
        1402 => x"83a50700",
        1403 => x"63860500",
        1404 => x"13050400",
        1405 => x"eff0dfbe",
        1406 => x"83254401",
        1407 => x"63860500",
        1408 => x"13050400",
        1409 => x"eff0dfbd",
        1410 => x"83254402",
        1411 => x"63860500",
        1412 => x"13050400",
        1413 => x"eff0dfbc",
        1414 => x"83258403",
        1415 => x"63860500",
        1416 => x"13050400",
        1417 => x"eff0dfbb",
        1418 => x"8325c403",
        1419 => x"63860500",
        1420 => x"13050400",
        1421 => x"eff0dfba",
        1422 => x"83250404",
        1423 => x"63860500",
        1424 => x"13050400",
        1425 => x"eff0dfb9",
        1426 => x"8325c405",
        1427 => x"63860500",
        1428 => x"13050400",
        1429 => x"eff0dfb8",
        1430 => x"83258405",
        1431 => x"63860500",
        1432 => x"13050400",
        1433 => x"eff0dfb7",
        1434 => x"83254403",
        1435 => x"63860500",
        1436 => x"13050400",
        1437 => x"eff0dfb6",
        1438 => x"83278401",
        1439 => x"638a0706",
        1440 => x"83278402",
        1441 => x"13050400",
        1442 => x"e7800700",
        1443 => x"83258404",
        1444 => x"63800506",
        1445 => x"13050400",
        1446 => x"03248101",
        1447 => x"8320c101",
        1448 => x"83244101",
        1449 => x"03290101",
        1450 => x"8329c100",
        1451 => x"13010102",
        1452 => x"6ff09feb",
        1453 => x"b3859500",
        1454 => x"83a50500",
        1455 => x"63900502",
        1456 => x"93844400",
        1457 => x"83274402",
        1458 => x"83a5c700",
        1459 => x"e39424ff",
        1460 => x"13050400",
        1461 => x"eff0dfb0",
        1462 => x"6ff0dff0",
        1463 => x"83a90500",
        1464 => x"13050400",
        1465 => x"eff0dfaf",
        1466 => x"93850900",
        1467 => x"6ff01ffd",
        1468 => x"8320c101",
        1469 => x"03248101",
        1470 => x"83244101",
        1471 => x"03290101",
        1472 => x"8329c100",
        1473 => x"13010102",
        1474 => x"67800000",
        1475 => x"67800000",
        1476 => x"57616974",
        1477 => x"2e2e2e2e",
        1478 => x"0d000000",
        1479 => x"35207365",
        1480 => x"636f6e64",
        1481 => x"7320656c",
        1482 => x"61707365",
        1483 => x"640d0a00",
        1484 => x"0d0a0d0a",
        1485 => x"496e7465",
        1486 => x"7276616c",
        1487 => x"20746573",
        1488 => x"74696e67",
        1489 => x"0d0a0000",
        1490 => x"436c6f63",
        1491 => x"6b732070",
        1492 => x"65722073",
        1493 => x"65636f6e",
        1494 => x"643a2025",
        1495 => x"640d0a00",
        1496 => x"256c750d",
        1497 => x"0a000000",
        1498 => x"232d302b",
        1499 => x"20000000",
        1500 => x"686c4c00",
        1501 => x"65666745",
        1502 => x"46470000",
        1503 => x"30313233",
        1504 => x"34353637",
        1505 => x"38394142",
        1506 => x"43444546",
        1507 => x"00000000",
        1508 => x"30313233",
        1509 => x"34353637",
        1510 => x"38396162",
        1511 => x"63646566",
        1512 => x"00000000",
        1513 => x"b40e0000",
        1514 => x"d40e0000",
        1515 => x"800e0000",
        1516 => x"800e0000",
        1517 => x"800e0000",
        1518 => x"800e0000",
        1519 => x"d40e0000",
        1520 => x"800e0000",
        1521 => x"800e0000",
        1522 => x"800e0000",
        1523 => x"800e0000",
        1524 => x"c0100000",
        1525 => x"2c0f0000",
        1526 => x"3c100000",
        1527 => x"800e0000",
        1528 => x"800e0000",
        1529 => x"08110000",
        1530 => x"800e0000",
        1531 => x"2c0f0000",
        1532 => x"800e0000",
        1533 => x"800e0000",
        1534 => x"48100000",
        1535 => x"00000020",
        1536 => x"00000000",
        1537 => x"00000000",
        1538 => x"00000000",
        1539 => x"00000000",
        1540 => x"00000000",
        1541 => x"00000000",
        1542 => x"00000000",
        1543 => x"00000000",
        1544 => x"00000000",
        1545 => x"00000000",
        1546 => x"00000000",
        1547 => x"00000000",
        1548 => x"00000000",
        1549 => x"00000000",
        1550 => x"00000000",
        1551 => x"00000000",
        1552 => x"00000000",
        1553 => x"00000000",
        1554 => x"00000000",
        1555 => x"00000000",
        1556 => x"00000000",
        1557 => x"00000000",
        1558 => x"00000000",
        1559 => x"00000000",
        1560 => x"00000020",
        others => (others => '0')
    );
end package processor_common_rom;
