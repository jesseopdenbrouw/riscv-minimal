-- srec2vhdl table generator
-- for input file main.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"93828206",
           6 => x"73905230",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef101000",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"93850532",
          21 => x"13050500",
          22 => x"ef10807b",
          23 => x"ef10d021",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10d001",
          29 => x"ef10501c",
          30 => x"6f000000",
          31 => x"37170000",
          32 => x"b70700f0",
          33 => x"13077745",
          34 => x"23a2e702",
          35 => x"13070004",
          36 => x"23a4e702",
          37 => x"67800000",
          38 => x"1375f50f",
          39 => x"b70700f0",
          40 => x"23a0a702",
          41 => x"370700f0",
          42 => x"8327c702",
          43 => x"93f70701",
          44 => x"e38c07fe",
          45 => x"67800000",
          46 => x"63060502",
          47 => x"83470500",
          48 => x"63820702",
          49 => x"370700f0",
          50 => x"13051500",
          51 => x"2320f702",
          52 => x"8327c702",
          53 => x"93f70701",
          54 => x"e38c07fe",
          55 => x"83470500",
          56 => x"e39407fe",
          57 => x"67800000",
          58 => x"370700f0",
          59 => x"8327c702",
          60 => x"93f74700",
          61 => x"e38c07fe",
          62 => x"03250702",
          63 => x"1375f50f",
          64 => x"67800000",
          65 => x"130101ff",
          66 => x"373e0000",
          67 => x"370700f0",
          68 => x"930e0500",
          69 => x"138ff5ff",
          70 => x"23268100",
          71 => x"13050000",
          72 => x"130ecef2",
          73 => x"13070702",
          74 => x"13035001",
          75 => x"93027000",
          76 => x"930fe005",
          77 => x"9305f007",
          78 => x"93082000",
          79 => x"13082001",
          80 => x"b7330000",
          81 => x"1306f007",
          82 => x"8327c700",
          83 => x"93f74700",
          84 => x"e38c07fe",
          85 => x"03240700",
          86 => x"9376f40f",
          87 => x"636ed302",
          88 => x"63fed802",
          89 => x"9387d6ff",
          90 => x"636af802",
          91 => x"93972700",
          92 => x"b307fe00",
          93 => x"83a70700",
          94 => x"67800700",
          95 => x"1305f5ff",
          96 => x"6308050c",
          97 => x"2320c700",
          98 => x"8327c700",
          99 => x"93f70701",
         100 => x"e38c07fe",
         101 => x"6ff09ffe",
         102 => x"638cb606",
         103 => x"635ae50d",
         104 => x"1374f40f",
         105 => x"930704fe",
         106 => x"93f7f70f",
         107 => x"e3eefff8",
         108 => x"b387ae00",
         109 => x"23808700",
         110 => x"13051500",
         111 => x"2320d700",
         112 => x"8327c700",
         113 => x"93f70701",
         114 => x"e38c07fe",
         115 => x"6ff0dff7",
         116 => x"b38eae00",
         117 => x"b7360000",
         118 => x"23800e00",
         119 => x"9307d000",
         120 => x"9386861a",
         121 => x"370700f0",
         122 => x"93861600",
         123 => x"2320f702",
         124 => x"8327c702",
         125 => x"93f70701",
         126 => x"e38c07fe",
         127 => x"83c70600",
         128 => x"e39407fe",
         129 => x"0324c100",
         130 => x"13010101",
         131 => x"67800000",
         132 => x"63040504",
         133 => x"2320b700",
         134 => x"8327c700",
         135 => x"93f70701",
         136 => x"e38c07fe",
         137 => x"1305f5ff",
         138 => x"6ff01ff2",
         139 => x"9307c003",
         140 => x"93868326",
         141 => x"93861600",
         142 => x"2320f700",
         143 => x"8327c700",
         144 => x"93f70701",
         145 => x"e38c07fe",
         146 => x"83c70600",
         147 => x"e39407fe",
         148 => x"13050000",
         149 => x"6ff05fef",
         150 => x"23205700",
         151 => x"8327c700",
         152 => x"93f70701",
         153 => x"e38c07fe",
         154 => x"13050000",
         155 => x"6ff0dfed",
         156 => x"23205700",
         157 => x"8327c700",
         158 => x"93f70701",
         159 => x"e38c07fe",
         160 => x"6ff09fec",
         161 => x"1375f50f",
         162 => x"b70700f0",
         163 => x"23a0a702",
         164 => x"370700f0",
         165 => x"8327c702",
         166 => x"93f70701",
         167 => x"e38c07fe",
         168 => x"13051000",
         169 => x"67800000",
         170 => x"370700f0",
         171 => x"8327c702",
         172 => x"93f74700",
         173 => x"e38c07fe",
         174 => x"03250702",
         175 => x"1375f50f",
         176 => x"67800000",
         177 => x"13050000",
         178 => x"67800000",
         179 => x"13050000",
         180 => x"67800000",
         181 => x"130101f8",
         182 => x"23221100",
         183 => x"23242100",
         184 => x"23263100",
         185 => x"23284100",
         186 => x"232a5100",
         187 => x"232c6100",
         188 => x"232e7100",
         189 => x"23208102",
         190 => x"23229102",
         191 => x"2324a102",
         192 => x"2326b102",
         193 => x"2328c102",
         194 => x"232ad102",
         195 => x"232ce102",
         196 => x"232ef102",
         197 => x"23200105",
         198 => x"23221105",
         199 => x"23242105",
         200 => x"23263105",
         201 => x"23284105",
         202 => x"232a5105",
         203 => x"232c6105",
         204 => x"232e7105",
         205 => x"23208107",
         206 => x"23229107",
         207 => x"2324a107",
         208 => x"2326b107",
         209 => x"2328c107",
         210 => x"232ad107",
         211 => x"232ce107",
         212 => x"232ef107",
         213 => x"f3272034",
         214 => x"37070080",
         215 => x"93067700",
         216 => x"6388d70c",
         217 => x"9306b000",
         218 => x"63e4f602",
         219 => x"13071000",
         220 => x"637cf70a",
         221 => x"63eaf60a",
         222 => x"37370000",
         223 => x"93972700",
         224 => x"130787f7",
         225 => x"b387e700",
         226 => x"83a70700",
         227 => x"67800700",
         228 => x"93061701",
         229 => x"6384d70a",
         230 => x"13072701",
         231 => x"6396e708",
         232 => x"ef000037",
         233 => x"03258102",
         234 => x"832fc107",
         235 => x"032f8107",
         236 => x"832e4107",
         237 => x"032e0107",
         238 => x"832dc106",
         239 => x"032d8106",
         240 => x"832c4106",
         241 => x"032c0106",
         242 => x"832bc105",
         243 => x"032b8105",
         244 => x"832a4105",
         245 => x"032a0105",
         246 => x"8329c104",
         247 => x"03298104",
         248 => x"83284104",
         249 => x"03280104",
         250 => x"8327c103",
         251 => x"03278103",
         252 => x"83264103",
         253 => x"03260103",
         254 => x"8325c102",
         255 => x"83244102",
         256 => x"03240102",
         257 => x"8323c101",
         258 => x"03238101",
         259 => x"83224101",
         260 => x"03220101",
         261 => x"8321c100",
         262 => x"03218100",
         263 => x"83204100",
         264 => x"13010108",
         265 => x"73002030",
         266 => x"03258102",
         267 => x"6ff0dff7",
         268 => x"ef00c029",
         269 => x"03258102",
         270 => x"6ff01ff7",
         271 => x"ef00c026",
         272 => x"03258102",
         273 => x"6ff05ff6",
         274 => x"9307600d",
         275 => x"6388f814",
         276 => x"9307900a",
         277 => x"6382f818",
         278 => x"63cc1703",
         279 => x"938878fc",
         280 => x"93074002",
         281 => x"63e81705",
         282 => x"b7370000",
         283 => x"938787fa",
         284 => x"93982800",
         285 => x"b388f800",
         286 => x"83a70800",
         287 => x"67800700",
         288 => x"13050100",
         289 => x"ef00c01b",
         290 => x"03258102",
         291 => x"6ff0dff1",
         292 => x"938808c0",
         293 => x"9307f000",
         294 => x"63ee1701",
         295 => x"b7370000",
         296 => x"9387c703",
         297 => x"93982800",
         298 => x"b388f800",
         299 => x"83a70800",
         300 => x"67800700",
         301 => x"ef10c057",
         302 => x"93078005",
         303 => x"2320f500",
         304 => x"9307f0ff",
         305 => x"13850700",
         306 => x"6ff01fee",
         307 => x"b7270000",
         308 => x"23a2f500",
         309 => x"93070000",
         310 => x"13850700",
         311 => x"6ff0dfec",
         312 => x"93070000",
         313 => x"13850700",
         314 => x"6ff01fec",
         315 => x"ef104054",
         316 => x"93079000",
         317 => x"2320f500",
         318 => x"9307f0ff",
         319 => x"13850700",
         320 => x"6ff09fea",
         321 => x"ef10c052",
         322 => x"9307f001",
         323 => x"2320f500",
         324 => x"9307f0ff",
         325 => x"13850700",
         326 => x"6ff01fe9",
         327 => x"ef104051",
         328 => x"9307d000",
         329 => x"2320f500",
         330 => x"9307f0ff",
         331 => x"13850700",
         332 => x"6ff09fe7",
         333 => x"ef10c04f",
         334 => x"93072000",
         335 => x"2320f500",
         336 => x"9307f0ff",
         337 => x"13850700",
         338 => x"6ff01fe6",
         339 => x"13090600",
         340 => x"13840500",
         341 => x"635cc000",
         342 => x"b384c500",
         343 => x"03450400",
         344 => x"13041400",
         345 => x"eff01fd2",
         346 => x"e39a84fe",
         347 => x"13050900",
         348 => x"6ff09fe3",
         349 => x"13090600",
         350 => x"13840500",
         351 => x"e358c0fe",
         352 => x"b384c500",
         353 => x"eff05fd2",
         354 => x"2300a400",
         355 => x"13041400",
         356 => x"e31a94fe",
         357 => x"13050900",
         358 => x"6ff01fe1",
         359 => x"63180500",
         360 => x"13858189",
         361 => x"13050500",
         362 => x"6ff01fe0",
         363 => x"b7870020",
         364 => x"93870700",
         365 => x"13070040",
         366 => x"b387e740",
         367 => x"e364f5fe",
         368 => x"ef100047",
         369 => x"9307c000",
         370 => x"2320f500",
         371 => x"1305f0ff",
         372 => x"13050500",
         373 => x"6ff05fdd",
         374 => x"13090000",
         375 => x"93040500",
         376 => x"13040900",
         377 => x"93090900",
         378 => x"93070900",
         379 => x"732410c8",
         380 => x"f32910c0",
         381 => x"f32710c8",
         382 => x"e31af4fe",
         383 => x"37460f00",
         384 => x"13060624",
         385 => x"93060000",
         386 => x"13850900",
         387 => x"93050400",
         388 => x"ef00d061",
         389 => x"37460f00",
         390 => x"23a4a400",
         391 => x"13060624",
         392 => x"93060000",
         393 => x"13850900",
         394 => x"93050400",
         395 => x"ef00101d",
         396 => x"23a0a400",
         397 => x"23a2b400",
         398 => x"13050900",
         399 => x"6ff0dfd6",
         400 => x"37350000",
         401 => x"130101ff",
         402 => x"13054527",
         403 => x"23261100",
         404 => x"23248100",
         405 => x"23229100",
         406 => x"23202101",
         407 => x"eff0dfa5",
         408 => x"73294034",
         409 => x"93040002",
         410 => x"37040080",
         411 => x"33758900",
         412 => x"3335a000",
         413 => x"13050503",
         414 => x"9384f4ff",
         415 => x"eff0dfa1",
         416 => x"13541400",
         417 => x"e39404fe",
         418 => x"03248100",
         419 => x"8320c100",
         420 => x"83244100",
         421 => x"03290100",
         422 => x"37350000",
         423 => x"1305851a",
         424 => x"13010101",
         425 => x"6ff05fa1",
         426 => x"b70700f0",
         427 => x"03a74708",
         428 => x"1377f7fe",
         429 => x"23a2e708",
         430 => x"03a74700",
         431 => x"13471700",
         432 => x"23a2e700",
         433 => x"67800000",
         434 => x"6f000000",
         435 => x"b70700f0",
         436 => x"83a5470f",
         437 => x"03a7070f",
         438 => x"b7860100",
         439 => x"1306f0ff",
         440 => x"9386066a",
         441 => x"23aec70e",
         442 => x"b306d700",
         443 => x"23acc70e",
         444 => x"33b7e600",
         445 => x"23acd70e",
         446 => x"3307b700",
         447 => x"23aee70e",
         448 => x"03a74700",
         449 => x"13472700",
         450 => x"23a2e700",
         451 => x"67800000",
         452 => x"370700f0",
         453 => x"8327c702",
         454 => x"93f74700",
         455 => x"638a0700",
         456 => x"83274700",
         457 => x"93c74700",
         458 => x"2322f700",
         459 => x"83270702",
         460 => x"67800000",
         461 => x"13030500",
         462 => x"138e0500",
         463 => x"93080000",
         464 => x"63dc0500",
         465 => x"b337a000",
         466 => x"330eb040",
         467 => x"330efe40",
         468 => x"3303a040",
         469 => x"9308f0ff",
         470 => x"63dc0600",
         471 => x"b337c000",
         472 => x"b306d040",
         473 => x"93c8f8ff",
         474 => x"b386f640",
         475 => x"3306c040",
         476 => x"13070600",
         477 => x"13080300",
         478 => x"93070e00",
         479 => x"639c0628",
         480 => x"b7350000",
         481 => x"9385c507",
         482 => x"6376ce0e",
         483 => x"b7060100",
         484 => x"6378d60c",
         485 => x"93360610",
         486 => x"93c61600",
         487 => x"93963600",
         488 => x"3355d600",
         489 => x"b385a500",
         490 => x"83c50500",
         491 => x"13050002",
         492 => x"b386d500",
         493 => x"b305d540",
         494 => x"630cd500",
         495 => x"b317be00",
         496 => x"b356d300",
         497 => x"3317b600",
         498 => x"b3e7f600",
         499 => x"3318b300",
         500 => x"93550701",
         501 => x"33deb702",
         502 => x"13160701",
         503 => x"13560601",
         504 => x"b3f7b702",
         505 => x"13050e00",
         506 => x"3303c603",
         507 => x"93960701",
         508 => x"93570801",
         509 => x"b3e7d700",
         510 => x"63fe6700",
         511 => x"b387e700",
         512 => x"1305feff",
         513 => x"63e8e700",
         514 => x"63f66700",
         515 => x"1305eeff",
         516 => x"b387e700",
         517 => x"b3876740",
         518 => x"33d3b702",
         519 => x"13180801",
         520 => x"13580801",
         521 => x"b3f7b702",
         522 => x"b3066602",
         523 => x"93970701",
         524 => x"3368f800",
         525 => x"93070300",
         526 => x"637cd800",
         527 => x"33080701",
         528 => x"9307f3ff",
         529 => x"6366e800",
         530 => x"6374d800",
         531 => x"9307e3ff",
         532 => x"13150501",
         533 => x"3365f500",
         534 => x"93050000",
         535 => x"6f00000e",
         536 => x"37050001",
         537 => x"93060001",
         538 => x"e36ca6f2",
         539 => x"93068001",
         540 => x"6ff01ff3",
         541 => x"63140600",
         542 => x"73001000",
         543 => x"b7070100",
         544 => x"637af60c",
         545 => x"93360610",
         546 => x"93c61600",
         547 => x"93963600",
         548 => x"b357d600",
         549 => x"b385f500",
         550 => x"83c70500",
         551 => x"b387d700",
         552 => x"93060002",
         553 => x"b385f640",
         554 => x"6390f60c",
         555 => x"b307ce40",
         556 => x"93051000",
         557 => x"13530701",
         558 => x"b3de6702",
         559 => x"13160701",
         560 => x"13560601",
         561 => x"93560801",
         562 => x"b3f76702",
         563 => x"13850e00",
         564 => x"330ed603",
         565 => x"93970701",
         566 => x"b3e7f600",
         567 => x"63fec701",
         568 => x"b387e700",
         569 => x"1385feff",
         570 => x"63e8e700",
         571 => x"63f6c701",
         572 => x"1385eeff",
         573 => x"b387e700",
         574 => x"b387c741",
         575 => x"33de6702",
         576 => x"13180801",
         577 => x"13580801",
         578 => x"b3f76702",
         579 => x"b306c603",
         580 => x"93970701",
         581 => x"3368f800",
         582 => x"93070e00",
         583 => x"637cd800",
         584 => x"33080701",
         585 => x"9307feff",
         586 => x"6366e800",
         587 => x"6374d800",
         588 => x"9307eeff",
         589 => x"13150501",
         590 => x"3365f500",
         591 => x"638a0800",
         592 => x"b337a000",
         593 => x"b305b040",
         594 => x"b385f540",
         595 => x"3305a040",
         596 => x"67800000",
         597 => x"b7070001",
         598 => x"93060001",
         599 => x"e36af6f2",
         600 => x"93068001",
         601 => x"6ff0dff2",
         602 => x"3317b600",
         603 => x"b356fe00",
         604 => x"13550701",
         605 => x"331ebe00",
         606 => x"b357f300",
         607 => x"b3e7c701",
         608 => x"33dea602",
         609 => x"13160701",
         610 => x"13560601",
         611 => x"3318b300",
         612 => x"b3f6a602",
         613 => x"3303c603",
         614 => x"93950601",
         615 => x"93d60701",
         616 => x"b3e6b600",
         617 => x"93050e00",
         618 => x"63fe6600",
         619 => x"b386e600",
         620 => x"9305feff",
         621 => x"63e8e600",
         622 => x"63f66600",
         623 => x"9305eeff",
         624 => x"b386e600",
         625 => x"b3866640",
         626 => x"33d3a602",
         627 => x"93970701",
         628 => x"93d70701",
         629 => x"b3f6a602",
         630 => x"33066602",
         631 => x"93960601",
         632 => x"b3e7d700",
         633 => x"93060300",
         634 => x"63fec700",
         635 => x"b387e700",
         636 => x"9306f3ff",
         637 => x"63e8e700",
         638 => x"63f6c700",
         639 => x"9306e3ff",
         640 => x"b387e700",
         641 => x"93950501",
         642 => x"b387c740",
         643 => x"b3e5d500",
         644 => x"6ff05fea",
         645 => x"6366de18",
         646 => x"b7070100",
         647 => x"63f4f604",
         648 => x"13b70610",
         649 => x"13471700",
         650 => x"13173700",
         651 => x"b7370000",
         652 => x"b3d5e600",
         653 => x"9387c707",
         654 => x"b387b700",
         655 => x"83c70700",
         656 => x"b387e700",
         657 => x"13070002",
         658 => x"b305f740",
         659 => x"6316f702",
         660 => x"13051000",
         661 => x"e3e4c6ef",
         662 => x"3335c300",
         663 => x"13451500",
         664 => x"6ff0dfed",
         665 => x"b7070001",
         666 => x"13070001",
         667 => x"e3e0f6fc",
         668 => x"13078001",
         669 => x"6ff09ffb",
         670 => x"3357f600",
         671 => x"b396b600",
         672 => x"b366d700",
         673 => x"3357fe00",
         674 => x"331ebe00",
         675 => x"b357f300",
         676 => x"b3e7c701",
         677 => x"13de0601",
         678 => x"335fc703",
         679 => x"13980601",
         680 => x"13580801",
         681 => x"3316b600",
         682 => x"3377c703",
         683 => x"b30ee803",
         684 => x"13150701",
         685 => x"13d70701",
         686 => x"3367a700",
         687 => x"13050f00",
         688 => x"637ed701",
         689 => x"3307d700",
         690 => x"1305ffff",
         691 => x"6368d700",
         692 => x"6376d701",
         693 => x"1305efff",
         694 => x"3307d700",
         695 => x"3307d741",
         696 => x"b35ec703",
         697 => x"93970701",
         698 => x"93d70701",
         699 => x"3377c703",
         700 => x"3308d803",
         701 => x"13170701",
         702 => x"b3e7e700",
         703 => x"13870e00",
         704 => x"63fe0701",
         705 => x"b387d700",
         706 => x"1387feff",
         707 => x"63e8d700",
         708 => x"63f60701",
         709 => x"1387eeff",
         710 => x"b387d700",
         711 => x"13150501",
         712 => x"b70e0100",
         713 => x"3365e500",
         714 => x"9386feff",
         715 => x"3377d500",
         716 => x"b3870741",
         717 => x"b376d600",
         718 => x"13580501",
         719 => x"13560601",
         720 => x"330ed702",
         721 => x"b306d802",
         722 => x"3307c702",
         723 => x"3308c802",
         724 => x"3306d700",
         725 => x"13570e01",
         726 => x"3307c700",
         727 => x"6374d700",
         728 => x"3308d801",
         729 => x"93560701",
         730 => x"b3860601",
         731 => x"63e6d702",
         732 => x"e394d7ce",
         733 => x"b7070100",
         734 => x"9387f7ff",
         735 => x"3377f700",
         736 => x"13170701",
         737 => x"337efe00",
         738 => x"3313b300",
         739 => x"3307c701",
         740 => x"93050000",
         741 => x"e374e3da",
         742 => x"1305f5ff",
         743 => x"6ff0dfcb",
         744 => x"93050000",
         745 => x"13050000",
         746 => x"6ff05fd9",
         747 => x"138e0500",
         748 => x"13080000",
         749 => x"63dc0500",
         750 => x"b337a000",
         751 => x"b305b040",
         752 => x"338ef540",
         753 => x"3305a040",
         754 => x"1308f0ff",
         755 => x"63da0600",
         756 => x"b337c000",
         757 => x"b306d040",
         758 => x"b386f640",
         759 => x"3306c040",
         760 => x"93080600",
         761 => x"93070500",
         762 => x"93050e00",
         763 => x"63940624",
         764 => x"37370000",
         765 => x"1307c707",
         766 => x"6376ce0e",
         767 => x"b7060100",
         768 => x"6378d60c",
         769 => x"93360610",
         770 => x"93c61600",
         771 => x"93963600",
         772 => x"3353d600",
         773 => x"33076700",
         774 => x"03470700",
         775 => x"3307d700",
         776 => x"93060002",
         777 => x"3383e640",
         778 => x"638ce600",
         779 => x"b3156e00",
         780 => x"3357e500",
         781 => x"b3186600",
         782 => x"b365b700",
         783 => x"b3176500",
         784 => x"93d60801",
         785 => x"33d7d502",
         786 => x"13950801",
         787 => x"13550501",
         788 => x"b3f5d502",
         789 => x"3307a702",
         790 => x"13960501",
         791 => x"93d50701",
         792 => x"b3e5c500",
         793 => x"63fae500",
         794 => x"b3851501",
         795 => x"63e61501",
         796 => x"63f4e500",
         797 => x"b3851501",
         798 => x"b385e540",
         799 => x"33d7d502",
         800 => x"93970701",
         801 => x"93d70701",
         802 => x"b3f5d502",
         803 => x"3307a702",
         804 => x"93950501",
         805 => x"b3e7b700",
         806 => x"63fae700",
         807 => x"b3871701",
         808 => x"63e61701",
         809 => x"63f4e700",
         810 => x"b3871701",
         811 => x"b387e740",
         812 => x"33d56700",
         813 => x"93050000",
         814 => x"630a0800",
         815 => x"b337a000",
         816 => x"b305b040",
         817 => x"b385f540",
         818 => x"3305a040",
         819 => x"67800000",
         820 => x"37030001",
         821 => x"93060001",
         822 => x"e36c66f2",
         823 => x"93068001",
         824 => x"6ff01ff3",
         825 => x"63140600",
         826 => x"73001000",
         827 => x"b7060100",
         828 => x"6372d60a",
         829 => x"93360610",
         830 => x"93c61600",
         831 => x"93963600",
         832 => x"b355d600",
         833 => x"3307b700",
         834 => x"03470700",
         835 => x"3307d700",
         836 => x"93060002",
         837 => x"3383e640",
         838 => x"6398e608",
         839 => x"3307ce40",
         840 => x"93d50801",
         841 => x"3356b702",
         842 => x"13950801",
         843 => x"13550501",
         844 => x"93d60701",
         845 => x"3377b702",
         846 => x"3306a602",
         847 => x"13170701",
         848 => x"33e7e600",
         849 => x"637ac700",
         850 => x"33071701",
         851 => x"63661701",
         852 => x"6374c700",
         853 => x"33071701",
         854 => x"3307c740",
         855 => x"b356b702",
         856 => x"93970701",
         857 => x"93d70701",
         858 => x"3377b702",
         859 => x"b386a602",
         860 => x"13170701",
         861 => x"b3e7e700",
         862 => x"63fad700",
         863 => x"b3871701",
         864 => x"63e61701",
         865 => x"63f4d700",
         866 => x"b3871701",
         867 => x"b387d740",
         868 => x"6ff01ff2",
         869 => x"b7050001",
         870 => x"93060001",
         871 => x"e362b6f6",
         872 => x"93068001",
         873 => x"6ff0dff5",
         874 => x"b3186600",
         875 => x"b356ee00",
         876 => x"b3156e00",
         877 => x"3357e500",
         878 => x"b3176500",
         879 => x"13d50801",
         880 => x"3367b700",
         881 => x"b3d5a602",
         882 => x"139e0801",
         883 => x"135e0e01",
         884 => x"b3f6a602",
         885 => x"b385c503",
         886 => x"13960601",
         887 => x"93560701",
         888 => x"b3e6c600",
         889 => x"63fab600",
         890 => x"b3861601",
         891 => x"63e61601",
         892 => x"63f4b600",
         893 => x"b3861601",
         894 => x"b386b640",
         895 => x"33d6a602",
         896 => x"13170701",
         897 => x"13570701",
         898 => x"b3f6a602",
         899 => x"3306c603",
         900 => x"93960601",
         901 => x"3367d700",
         902 => x"637ac700",
         903 => x"33071701",
         904 => x"63661701",
         905 => x"6374c700",
         906 => x"33071701",
         907 => x"3307c740",
         908 => x"6ff01fef",
         909 => x"e362dee8",
         910 => x"37070100",
         911 => x"63fce604",
         912 => x"13b70610",
         913 => x"13471700",
         914 => x"13173700",
         915 => x"b7380000",
         916 => x"33d3e600",
         917 => x"9388c807",
         918 => x"b3886800",
         919 => x"03c30800",
         920 => x"3303e300",
         921 => x"13070002",
         922 => x"b3086740",
         923 => x"631e6702",
         924 => x"63e4c601",
         925 => x"636cc500",
         926 => x"3306c540",
         927 => x"b306de40",
         928 => x"b335c500",
         929 => x"b385b640",
         930 => x"93070600",
         931 => x"13850700",
         932 => x"6ff09fe2",
         933 => x"b7080001",
         934 => x"13070001",
         935 => x"e3e816fb",
         936 => x"13078001",
         937 => x"6ff09ffa",
         938 => x"b3576600",
         939 => x"b3961601",
         940 => x"b3e6d700",
         941 => x"33576e00",
         942 => x"93de0601",
         943 => x"b35fd703",
         944 => x"b3151e01",
         945 => x"139e0601",
         946 => x"135e0e01",
         947 => x"b3576500",
         948 => x"b3e5b700",
         949 => x"93d70501",
         950 => x"33161601",
         951 => x"33151501",
         952 => x"3377d703",
         953 => x"330ffe03",
         954 => x"13170701",
         955 => x"b3e7e700",
         956 => x"13870f00",
         957 => x"63fee701",
         958 => x"b387d700",
         959 => x"1387ffff",
         960 => x"63e8d700",
         961 => x"63f6e701",
         962 => x"1387efff",
         963 => x"b387d700",
         964 => x"b387e741",
         965 => x"33dfd703",
         966 => x"93950501",
         967 => x"93d50501",
         968 => x"b3f7d703",
         969 => x"330eee03",
         970 => x"93970701",
         971 => x"b3e5f500",
         972 => x"93070f00",
         973 => x"63fec501",
         974 => x"b385d500",
         975 => x"9307ffff",
         976 => x"63e8d500",
         977 => x"63f6c501",
         978 => x"9307efff",
         979 => x"b385d500",
         980 => x"13170701",
         981 => x"b70f0100",
         982 => x"3367f700",
         983 => x"b385c541",
         984 => x"138effff",
         985 => x"b377c701",
         986 => x"935e0601",
         987 => x"13570701",
         988 => x"337ec601",
         989 => x"338fc703",
         990 => x"330ec703",
         991 => x"b387d703",
         992 => x"3307d703",
         993 => x"b38ec701",
         994 => x"93570f01",
         995 => x"b387d701",
         996 => x"63f4c701",
         997 => x"3307f701",
         998 => x"13de0701",
         999 => x"3307ee00",
        1000 => x"370e0100",
        1001 => x"130efeff",
        1002 => x"b3f7c701",
        1003 => x"93970701",
        1004 => x"337fcf01",
        1005 => x"b387e701",
        1006 => x"63e6e500",
        1007 => x"639ee500",
        1008 => x"637cf500",
        1009 => x"3386c740",
        1010 => x"b3b7c700",
        1011 => x"b387d700",
        1012 => x"3307f740",
        1013 => x"93070600",
        1014 => x"b307f540",
        1015 => x"3335f500",
        1016 => x"b385e540",
        1017 => x"b385a540",
        1018 => x"33936500",
        1019 => x"b3d71701",
        1020 => x"3365f300",
        1021 => x"b3d51501",
        1022 => x"6ff01fcc",
        1023 => x"13030500",
        1024 => x"93880500",
        1025 => x"13070600",
        1026 => x"13080500",
        1027 => x"93870500",
        1028 => x"63920628",
        1029 => x"b7350000",
        1030 => x"9385c507",
        1031 => x"63f6c80e",
        1032 => x"b7060100",
        1033 => x"6378d60c",
        1034 => x"93360610",
        1035 => x"93c61600",
        1036 => x"93963600",
        1037 => x"3355d600",
        1038 => x"b385a500",
        1039 => x"83c50500",
        1040 => x"13050002",
        1041 => x"b386d500",
        1042 => x"b305d540",
        1043 => x"630cd500",
        1044 => x"b397b800",
        1045 => x"b356d300",
        1046 => x"3317b600",
        1047 => x"b3e7f600",
        1048 => x"3318b300",
        1049 => x"93550701",
        1050 => x"33d3b702",
        1051 => x"13160701",
        1052 => x"13560601",
        1053 => x"b3f7b702",
        1054 => x"13050300",
        1055 => x"b3086602",
        1056 => x"93960701",
        1057 => x"93570801",
        1058 => x"b3e7d700",
        1059 => x"63fe1701",
        1060 => x"b387e700",
        1061 => x"1305f3ff",
        1062 => x"63e8e700",
        1063 => x"63f61701",
        1064 => x"1305e3ff",
        1065 => x"b387e700",
        1066 => x"b3871741",
        1067 => x"b3d8b702",
        1068 => x"13180801",
        1069 => x"13580801",
        1070 => x"b3f7b702",
        1071 => x"b3061603",
        1072 => x"93970701",
        1073 => x"3368f800",
        1074 => x"93870800",
        1075 => x"637cd800",
        1076 => x"33080701",
        1077 => x"9387f8ff",
        1078 => x"6366e800",
        1079 => x"6374d800",
        1080 => x"9387e8ff",
        1081 => x"13150501",
        1082 => x"3365f500",
        1083 => x"93050000",
        1084 => x"67800000",
        1085 => x"37050001",
        1086 => x"93060001",
        1087 => x"e36ca6f2",
        1088 => x"93068001",
        1089 => x"6ff01ff3",
        1090 => x"63140600",
        1091 => x"73001000",
        1092 => x"b7070100",
        1093 => x"6370f60c",
        1094 => x"93360610",
        1095 => x"93c61600",
        1096 => x"93963600",
        1097 => x"b357d600",
        1098 => x"b385f500",
        1099 => x"83c70500",
        1100 => x"b387d700",
        1101 => x"93060002",
        1102 => x"b385f640",
        1103 => x"6396f60a",
        1104 => x"b387c840",
        1105 => x"93051000",
        1106 => x"93580701",
        1107 => x"33de1703",
        1108 => x"13160701",
        1109 => x"13560601",
        1110 => x"93560801",
        1111 => x"b3f71703",
        1112 => x"13050e00",
        1113 => x"3303c603",
        1114 => x"93970701",
        1115 => x"b3e7f600",
        1116 => x"63fe6700",
        1117 => x"b387e700",
        1118 => x"1305feff",
        1119 => x"63e8e700",
        1120 => x"63f66700",
        1121 => x"1305eeff",
        1122 => x"b387e700",
        1123 => x"b3876740",
        1124 => x"33d31703",
        1125 => x"13180801",
        1126 => x"13580801",
        1127 => x"b3f71703",
        1128 => x"b3066602",
        1129 => x"93970701",
        1130 => x"3368f800",
        1131 => x"93070300",
        1132 => x"637cd800",
        1133 => x"33080701",
        1134 => x"9307f3ff",
        1135 => x"6366e800",
        1136 => x"6374d800",
        1137 => x"9307e3ff",
        1138 => x"13150501",
        1139 => x"3365f500",
        1140 => x"67800000",
        1141 => x"b7070001",
        1142 => x"93060001",
        1143 => x"e364f6f4",
        1144 => x"93068001",
        1145 => x"6ff01ff4",
        1146 => x"3317b600",
        1147 => x"b3d6f800",
        1148 => x"13550701",
        1149 => x"b357f300",
        1150 => x"3318b300",
        1151 => x"33d3a602",
        1152 => x"13160701",
        1153 => x"b398b800",
        1154 => x"13560601",
        1155 => x"b3e71701",
        1156 => x"b3f6a602",
        1157 => x"b3086602",
        1158 => x"93950601",
        1159 => x"93d60701",
        1160 => x"b3e6b600",
        1161 => x"93050300",
        1162 => x"63fe1601",
        1163 => x"b386e600",
        1164 => x"9305f3ff",
        1165 => x"63e8e600",
        1166 => x"63f61601",
        1167 => x"9305e3ff",
        1168 => x"b386e600",
        1169 => x"b3861641",
        1170 => x"b3d8a602",
        1171 => x"93970701",
        1172 => x"93d70701",
        1173 => x"b3f6a602",
        1174 => x"33061603",
        1175 => x"93960601",
        1176 => x"b3e7d700",
        1177 => x"93860800",
        1178 => x"63fec700",
        1179 => x"b387e700",
        1180 => x"9386f8ff",
        1181 => x"63e8e700",
        1182 => x"63f6c700",
        1183 => x"9386e8ff",
        1184 => x"b387e700",
        1185 => x"93950501",
        1186 => x"b387c740",
        1187 => x"b3e5d500",
        1188 => x"6ff09feb",
        1189 => x"63e6d518",
        1190 => x"b7070100",
        1191 => x"63f4f604",
        1192 => x"13b70610",
        1193 => x"13471700",
        1194 => x"13173700",
        1195 => x"b7370000",
        1196 => x"b3d5e600",
        1197 => x"9387c707",
        1198 => x"b387b700",
        1199 => x"83c70700",
        1200 => x"b387e700",
        1201 => x"13070002",
        1202 => x"b305f740",
        1203 => x"6316f702",
        1204 => x"13051000",
        1205 => x"e3ee16e1",
        1206 => x"3335c300",
        1207 => x"13451500",
        1208 => x"67800000",
        1209 => x"b7070001",
        1210 => x"13070001",
        1211 => x"e3e0f6fc",
        1212 => x"13078001",
        1213 => x"6ff09ffb",
        1214 => x"3357f600",
        1215 => x"b396b600",
        1216 => x"b366d700",
        1217 => x"33d7f800",
        1218 => x"b398b800",
        1219 => x"b357f300",
        1220 => x"b3e71701",
        1221 => x"93d80601",
        1222 => x"b35e1703",
        1223 => x"13980601",
        1224 => x"13580801",
        1225 => x"3316b600",
        1226 => x"33771703",
        1227 => x"330ed803",
        1228 => x"13150701",
        1229 => x"13d70701",
        1230 => x"3367a700",
        1231 => x"13850e00",
        1232 => x"637ec701",
        1233 => x"3307d700",
        1234 => x"1385feff",
        1235 => x"6368d700",
        1236 => x"6376c701",
        1237 => x"1385eeff",
        1238 => x"3307d700",
        1239 => x"3307c741",
        1240 => x"335e1703",
        1241 => x"93970701",
        1242 => x"93d70701",
        1243 => x"33771703",
        1244 => x"3308c803",
        1245 => x"13170701",
        1246 => x"b3e7e700",
        1247 => x"13070e00",
        1248 => x"63fe0701",
        1249 => x"b387d700",
        1250 => x"1307feff",
        1251 => x"63e8d700",
        1252 => x"63f60701",
        1253 => x"1307eeff",
        1254 => x"b387d700",
        1255 => x"13150501",
        1256 => x"370e0100",
        1257 => x"3365e500",
        1258 => x"9306feff",
        1259 => x"3377d500",
        1260 => x"b3870741",
        1261 => x"b376d600",
        1262 => x"13580501",
        1263 => x"13560601",
        1264 => x"b308d702",
        1265 => x"b306d802",
        1266 => x"3307c702",
        1267 => x"3308c802",
        1268 => x"3306d700",
        1269 => x"13d70801",
        1270 => x"3307c700",
        1271 => x"6374d700",
        1272 => x"3308c801",
        1273 => x"93560701",
        1274 => x"b3860601",
        1275 => x"63e6d702",
        1276 => x"e39ed7ce",
        1277 => x"b7070100",
        1278 => x"9387f7ff",
        1279 => x"3377f700",
        1280 => x"13170701",
        1281 => x"b3f8f800",
        1282 => x"3313b300",
        1283 => x"33071701",
        1284 => x"93050000",
        1285 => x"e37ee3cc",
        1286 => x"1305f5ff",
        1287 => x"6ff01fcd",
        1288 => x"93050000",
        1289 => x"13050000",
        1290 => x"67800000",
        1291 => x"13080600",
        1292 => x"93070500",
        1293 => x"13870500",
        1294 => x"63960620",
        1295 => x"b7380000",
        1296 => x"9388c807",
        1297 => x"63fcc50c",
        1298 => x"b7060100",
        1299 => x"637ed60a",
        1300 => x"93360610",
        1301 => x"93c61600",
        1302 => x"93963600",
        1303 => x"3353d600",
        1304 => x"b3886800",
        1305 => x"83c80800",
        1306 => x"13030002",
        1307 => x"b386d800",
        1308 => x"b308d340",
        1309 => x"630cd300",
        1310 => x"33971501",
        1311 => x"b356d500",
        1312 => x"33181601",
        1313 => x"33e7e600",
        1314 => x"b3171501",
        1315 => x"13560801",
        1316 => x"b356c702",
        1317 => x"13150801",
        1318 => x"13550501",
        1319 => x"3377c702",
        1320 => x"b386a602",
        1321 => x"93150701",
        1322 => x"13d70701",
        1323 => x"3367b700",
        1324 => x"637ad700",
        1325 => x"33070701",
        1326 => x"63660701",
        1327 => x"6374d700",
        1328 => x"33070701",
        1329 => x"3307d740",
        1330 => x"b356c702",
        1331 => x"3377c702",
        1332 => x"b386a602",
        1333 => x"93970701",
        1334 => x"13170701",
        1335 => x"93d70701",
        1336 => x"b3e7e700",
        1337 => x"63fad700",
        1338 => x"b3870701",
        1339 => x"63e60701",
        1340 => x"63f4d700",
        1341 => x"b3870701",
        1342 => x"b387d740",
        1343 => x"33d51701",
        1344 => x"93050000",
        1345 => x"67800000",
        1346 => x"37030001",
        1347 => x"93060001",
        1348 => x"e36666f4",
        1349 => x"93068001",
        1350 => x"6ff05ff4",
        1351 => x"63140600",
        1352 => x"73001000",
        1353 => x"37070100",
        1354 => x"637ee606",
        1355 => x"93360610",
        1356 => x"93c61600",
        1357 => x"93963600",
        1358 => x"3357d600",
        1359 => x"b388e800",
        1360 => x"03c70800",
        1361 => x"3307d700",
        1362 => x"93060002",
        1363 => x"b388e640",
        1364 => x"6394e606",
        1365 => x"3387c540",
        1366 => x"93550801",
        1367 => x"3356b702",
        1368 => x"13150801",
        1369 => x"13550501",
        1370 => x"93d60701",
        1371 => x"3377b702",
        1372 => x"3306a602",
        1373 => x"13170701",
        1374 => x"33e7e600",
        1375 => x"637ac700",
        1376 => x"33070701",
        1377 => x"63660701",
        1378 => x"6374c700",
        1379 => x"33070701",
        1380 => x"3307c740",
        1381 => x"b356b702",
        1382 => x"3377b702",
        1383 => x"b386a602",
        1384 => x"6ff05ff3",
        1385 => x"37070001",
        1386 => x"93060001",
        1387 => x"e366e6f8",
        1388 => x"93068001",
        1389 => x"6ff05ff8",
        1390 => x"33181601",
        1391 => x"b3d6e500",
        1392 => x"b3171501",
        1393 => x"b3951501",
        1394 => x"3357e500",
        1395 => x"13550801",
        1396 => x"3367b700",
        1397 => x"b3d5a602",
        1398 => x"13130801",
        1399 => x"13530301",
        1400 => x"b3f6a602",
        1401 => x"b3856502",
        1402 => x"13960601",
        1403 => x"93560701",
        1404 => x"b3e6c600",
        1405 => x"63fab600",
        1406 => x"b3860601",
        1407 => x"63e60601",
        1408 => x"63f4b600",
        1409 => x"b3860601",
        1410 => x"b386b640",
        1411 => x"33d6a602",
        1412 => x"13170701",
        1413 => x"13570701",
        1414 => x"b3f6a602",
        1415 => x"33066602",
        1416 => x"93960601",
        1417 => x"3367d700",
        1418 => x"637ac700",
        1419 => x"33070701",
        1420 => x"63660701",
        1421 => x"6374c700",
        1422 => x"33070701",
        1423 => x"3307c740",
        1424 => x"6ff09ff1",
        1425 => x"63e4d51c",
        1426 => x"37080100",
        1427 => x"63fe0605",
        1428 => x"13b80610",
        1429 => x"13481800",
        1430 => x"13183800",
        1431 => x"b7380000",
        1432 => x"33d30601",
        1433 => x"9388c807",
        1434 => x"b3886800",
        1435 => x"83c80800",
        1436 => x"13030002",
        1437 => x"b3880801",
        1438 => x"33081341",
        1439 => x"63101305",
        1440 => x"63e4b600",
        1441 => x"636cc500",
        1442 => x"3306c540",
        1443 => x"b386d540",
        1444 => x"3337c500",
        1445 => x"3387e640",
        1446 => x"93070600",
        1447 => x"13850700",
        1448 => x"93050700",
        1449 => x"67800000",
        1450 => x"b7080001",
        1451 => x"13080001",
        1452 => x"e3e616fb",
        1453 => x"13088001",
        1454 => x"6ff05ffa",
        1455 => x"b3960601",
        1456 => x"33531601",
        1457 => x"3363d300",
        1458 => x"135e0301",
        1459 => x"b3d61501",
        1460 => x"33dfc603",
        1461 => x"13170301",
        1462 => x"13570701",
        1463 => x"b3970501",
        1464 => x"b3551501",
        1465 => x"b3e5f500",
        1466 => x"93d70501",
        1467 => x"33160601",
        1468 => x"33150501",
        1469 => x"b3f6c603",
        1470 => x"b30ee703",
        1471 => x"93960601",
        1472 => x"b3e7d700",
        1473 => x"93060f00",
        1474 => x"63fed701",
        1475 => x"b3876700",
        1476 => x"9306ffff",
        1477 => x"63e86700",
        1478 => x"63f6d701",
        1479 => x"9306efff",
        1480 => x"b3876700",
        1481 => x"b387d741",
        1482 => x"b3dec703",
        1483 => x"93950501",
        1484 => x"93d50501",
        1485 => x"b3f7c703",
        1486 => x"3307d703",
        1487 => x"93970701",
        1488 => x"b3e5f500",
        1489 => x"93870e00",
        1490 => x"63fee500",
        1491 => x"b3856500",
        1492 => x"9387feff",
        1493 => x"63e86500",
        1494 => x"63f6e500",
        1495 => x"9387eeff",
        1496 => x"b3856500",
        1497 => x"93960601",
        1498 => x"370f0100",
        1499 => x"b3e6f600",
        1500 => x"9307ffff",
        1501 => x"135e0601",
        1502 => x"b385e540",
        1503 => x"33f7f600",
        1504 => x"93d60601",
        1505 => x"b377f600",
        1506 => x"b30ef702",
        1507 => x"b387f602",
        1508 => x"3307c703",
        1509 => x"b386c603",
        1510 => x"330ef700",
        1511 => x"13d70e01",
        1512 => x"3307c701",
        1513 => x"6374f700",
        1514 => x"b386e601",
        1515 => x"93570701",
        1516 => x"b387d700",
        1517 => x"b7060100",
        1518 => x"9386f6ff",
        1519 => x"3377d700",
        1520 => x"13170701",
        1521 => x"b3fede00",
        1522 => x"3307d701",
        1523 => x"63e6f500",
        1524 => x"639ef500",
        1525 => x"637ce500",
        1526 => x"3306c740",
        1527 => x"3337c700",
        1528 => x"33076700",
        1529 => x"b387e740",
        1530 => x"13070600",
        1531 => x"3307e540",
        1532 => x"3335e500",
        1533 => x"b385f540",
        1534 => x"b385a540",
        1535 => x"b3981501",
        1536 => x"33570701",
        1537 => x"33e5e800",
        1538 => x"b3d50501",
        1539 => x"67800000",
        1540 => x"13030500",
        1541 => x"630e0600",
        1542 => x"83830500",
        1543 => x"23007300",
        1544 => x"1306f6ff",
        1545 => x"13031300",
        1546 => x"93851500",
        1547 => x"e31606fe",
        1548 => x"67800000",
        1549 => x"13030500",
        1550 => x"630a0600",
        1551 => x"2300b300",
        1552 => x"1306f6ff",
        1553 => x"13031300",
        1554 => x"e31a06fe",
        1555 => x"67800000",
        1556 => x"630c0602",
        1557 => x"13030500",
        1558 => x"93061000",
        1559 => x"636ab500",
        1560 => x"9306f0ff",
        1561 => x"1307f6ff",
        1562 => x"3303e300",
        1563 => x"b385e500",
        1564 => x"83830500",
        1565 => x"23007300",
        1566 => x"1306f6ff",
        1567 => x"3303d300",
        1568 => x"b385d500",
        1569 => x"e31606fe",
        1570 => x"67800000",
        1571 => x"130101f9",
        1572 => x"23248106",
        1573 => x"232e3105",
        1574 => x"23261106",
        1575 => x"23229106",
        1576 => x"23202107",
        1577 => x"232c4105",
        1578 => x"232a5105",
        1579 => x"23286105",
        1580 => x"23267105",
        1581 => x"23248105",
        1582 => x"93090500",
        1583 => x"13840500",
        1584 => x"232c0100",
        1585 => x"232e0100",
        1586 => x"23200102",
        1587 => x"23220102",
        1588 => x"23240102",
        1589 => x"23260102",
        1590 => x"23280102",
        1591 => x"232a0102",
        1592 => x"232c0102",
        1593 => x"232e0102",
        1594 => x"97f2ffff",
        1595 => x"9382c29e",
        1596 => x"73905230",
        1597 => x"b7220000",
        1598 => x"93828280",
        1599 => x"73900230",
        1600 => x"efe0cff7",
        1601 => x"b7877d01",
        1602 => x"370700f0",
        1603 => x"9387f783",
        1604 => x"2326f708",
        1605 => x"37390000",
        1606 => x"93071001",
        1607 => x"2320f708",
        1608 => x"1305891a",
        1609 => x"efe04ff9",
        1610 => x"63543003",
        1611 => x"9384f9ff",
        1612 => x"9309f0ff",
        1613 => x"03250400",
        1614 => x"9384f4ff",
        1615 => x"13044400",
        1616 => x"efe08ff7",
        1617 => x"1305891a",
        1618 => x"efe00ff7",
        1619 => x"e39434ff",
        1620 => x"37350000",
        1621 => x"1305c517",
        1622 => x"371a0000",
        1623 => x"efe0cff5",
        1624 => x"13040000",
        1625 => x"373c0000",
        1626 => x"130a0ae1",
        1627 => x"930a0000",
        1628 => x"930b0019",
        1629 => x"93050000",
        1630 => x"13058100",
        1631 => x"ef00c026",
        1632 => x"13041400",
        1633 => x"63020502",
        1634 => x"e31674ff",
        1635 => x"73001000",
        1636 => x"93050000",
        1637 => x"13058100",
        1638 => x"13040000",
        1639 => x"ef00c024",
        1640 => x"13041400",
        1641 => x"e31205fe",
        1642 => x"83248100",
        1643 => x"032bc100",
        1644 => x"1306c003",
        1645 => x"93060000",
        1646 => x"13850400",
        1647 => x"93050b00",
        1648 => x"eff0cf9e",
        1649 => x"93090500",
        1650 => x"1306c003",
        1651 => x"93060000",
        1652 => x"13850400",
        1653 => x"93050b00",
        1654 => x"efe0dfd5",
        1655 => x"1306c003",
        1656 => x"93060000",
        1657 => x"eff08f9c",
        1658 => x"13060a00",
        1659 => x"93860a00",
        1660 => x"13090500",
        1661 => x"93050b00",
        1662 => x"13850400",
        1663 => x"efe09fd3",
        1664 => x"83260101",
        1665 => x"13070500",
        1666 => x"13880900",
        1667 => x"93070900",
        1668 => x"13860400",
        1669 => x"9305cc1a",
        1670 => x"13058101",
        1671 => x"ef00c015",
        1672 => x"13058101",
        1673 => x"efe04fe9",
        1674 => x"e31674f5",
        1675 => x"6ff01ff6",
        1676 => x"03a5c187",
        1677 => x"67800000",
        1678 => x"130101ff",
        1679 => x"23248100",
        1680 => x"23261100",
        1681 => x"93070000",
        1682 => x"13040500",
        1683 => x"63880700",
        1684 => x"93050000",
        1685 => x"97000000",
        1686 => x"e7000000",
        1687 => x"b7370000",
        1688 => x"03a5c731",
        1689 => x"83278502",
        1690 => x"63840700",
        1691 => x"e7800700",
        1692 => x"13050400",
        1693 => x"ef108033",
        1694 => x"130101ff",
        1695 => x"23248100",
        1696 => x"23229100",
        1697 => x"37340000",
        1698 => x"b7340000",
        1699 => x"93870432",
        1700 => x"13040432",
        1701 => x"3304f440",
        1702 => x"23202101",
        1703 => x"23261100",
        1704 => x"13542440",
        1705 => x"93840432",
        1706 => x"13090000",
        1707 => x"63108904",
        1708 => x"b7340000",
        1709 => x"37340000",
        1710 => x"93870432",
        1711 => x"13040432",
        1712 => x"3304f440",
        1713 => x"13542440",
        1714 => x"93840432",
        1715 => x"13090000",
        1716 => x"63188902",
        1717 => x"8320c100",
        1718 => x"03248100",
        1719 => x"83244100",
        1720 => x"03290100",
        1721 => x"13010101",
        1722 => x"67800000",
        1723 => x"83a70400",
        1724 => x"13091900",
        1725 => x"93844400",
        1726 => x"e7800700",
        1727 => x"6ff01ffb",
        1728 => x"83a70400",
        1729 => x"13091900",
        1730 => x"93844400",
        1731 => x"e7800700",
        1732 => x"6ff01ffc",
        1733 => x"130101f6",
        1734 => x"232af108",
        1735 => x"b7070080",
        1736 => x"93c7f7ff",
        1737 => x"232ef100",
        1738 => x"2328f100",
        1739 => x"b707ffff",
        1740 => x"2326d108",
        1741 => x"2324b100",
        1742 => x"232cb100",
        1743 => x"93878720",
        1744 => x"9306c108",
        1745 => x"93058100",
        1746 => x"232e1106",
        1747 => x"232af100",
        1748 => x"2328e108",
        1749 => x"232c0109",
        1750 => x"232e1109",
        1751 => x"2322d100",
        1752 => x"ef004041",
        1753 => x"83278100",
        1754 => x"23800700",
        1755 => x"8320c107",
        1756 => x"1301010a",
        1757 => x"67800000",
        1758 => x"130101f6",
        1759 => x"232af108",
        1760 => x"b7070080",
        1761 => x"93c7f7ff",
        1762 => x"232ef100",
        1763 => x"2328f100",
        1764 => x"b707ffff",
        1765 => x"93878720",
        1766 => x"232af100",
        1767 => x"2324a100",
        1768 => x"232ca100",
        1769 => x"03a5c187",
        1770 => x"2324c108",
        1771 => x"2326d108",
        1772 => x"13860500",
        1773 => x"93068108",
        1774 => x"93058100",
        1775 => x"232e1106",
        1776 => x"2328e108",
        1777 => x"232c0109",
        1778 => x"232e1109",
        1779 => x"2322d100",
        1780 => x"ef00403a",
        1781 => x"83278100",
        1782 => x"23800700",
        1783 => x"8320c107",
        1784 => x"1301010a",
        1785 => x"67800000",
        1786 => x"13860500",
        1787 => x"93050500",
        1788 => x"03a5c187",
        1789 => x"6f004000",
        1790 => x"130101ff",
        1791 => x"23248100",
        1792 => x"23229100",
        1793 => x"13040500",
        1794 => x"13850500",
        1795 => x"93050600",
        1796 => x"23261100",
        1797 => x"23a20188",
        1798 => x"ef10401c",
        1799 => x"9307f0ff",
        1800 => x"6318f500",
        1801 => x"83a74188",
        1802 => x"63840700",
        1803 => x"2320f400",
        1804 => x"8320c100",
        1805 => x"03248100",
        1806 => x"83244100",
        1807 => x"13010101",
        1808 => x"67800000",
        1809 => x"130101fe",
        1810 => x"23282101",
        1811 => x"03a98500",
        1812 => x"232c8100",
        1813 => x"23263101",
        1814 => x"23244101",
        1815 => x"23225101",
        1816 => x"232e1100",
        1817 => x"232a9100",
        1818 => x"23206101",
        1819 => x"83aa0500",
        1820 => x"13840500",
        1821 => x"130a0600",
        1822 => x"93890600",
        1823 => x"63ec2609",
        1824 => x"83d7c500",
        1825 => x"13f70748",
        1826 => x"63040708",
        1827 => x"03274401",
        1828 => x"93043000",
        1829 => x"83a50501",
        1830 => x"b384e402",
        1831 => x"13072000",
        1832 => x"b38aba40",
        1833 => x"130b0500",
        1834 => x"b3c4e402",
        1835 => x"13871600",
        1836 => x"33075701",
        1837 => x"63f4e400",
        1838 => x"93040700",
        1839 => x"93f70740",
        1840 => x"6386070a",
        1841 => x"93850400",
        1842 => x"13050b00",
        1843 => x"ef001065",
        1844 => x"13090500",
        1845 => x"630c050a",
        1846 => x"83250401",
        1847 => x"13860a00",
        1848 => x"eff01fb3",
        1849 => x"8357c400",
        1850 => x"93f7f7b7",
        1851 => x"93e70708",
        1852 => x"2316f400",
        1853 => x"23282401",
        1854 => x"232a9400",
        1855 => x"33095901",
        1856 => x"b3845441",
        1857 => x"23202401",
        1858 => x"23249400",
        1859 => x"13890900",
        1860 => x"63f42901",
        1861 => x"13890900",
        1862 => x"03250400",
        1863 => x"13060900",
        1864 => x"93050a00",
        1865 => x"eff0dfb2",
        1866 => x"83278400",
        1867 => x"13050000",
        1868 => x"b3872741",
        1869 => x"2324f400",
        1870 => x"83270400",
        1871 => x"b3872701",
        1872 => x"2320f400",
        1873 => x"8320c101",
        1874 => x"03248101",
        1875 => x"83244101",
        1876 => x"03290101",
        1877 => x"8329c100",
        1878 => x"032a8100",
        1879 => x"832a4100",
        1880 => x"032b0100",
        1881 => x"13010102",
        1882 => x"67800000",
        1883 => x"13860400",
        1884 => x"13050b00",
        1885 => x"ef00906f",
        1886 => x"13090500",
        1887 => x"e31c05f6",
        1888 => x"83250401",
        1889 => x"13050b00",
        1890 => x"ef00d049",
        1891 => x"9307c000",
        1892 => x"2320fb00",
        1893 => x"8357c400",
        1894 => x"1305f0ff",
        1895 => x"93e70704",
        1896 => x"2316f400",
        1897 => x"6ff01ffa",
        1898 => x"83278600",
        1899 => x"130101fd",
        1900 => x"232e3101",
        1901 => x"23286101",
        1902 => x"23261102",
        1903 => x"23248102",
        1904 => x"23229102",
        1905 => x"23202103",
        1906 => x"232c4101",
        1907 => x"232a5101",
        1908 => x"23267101",
        1909 => x"23248101",
        1910 => x"23229101",
        1911 => x"2320a101",
        1912 => x"032b0600",
        1913 => x"93090600",
        1914 => x"63980712",
        1915 => x"13050000",
        1916 => x"8320c102",
        1917 => x"03248102",
        1918 => x"23a20900",
        1919 => x"83244102",
        1920 => x"03290102",
        1921 => x"8329c101",
        1922 => x"032a8101",
        1923 => x"832a4101",
        1924 => x"032b0101",
        1925 => x"832bc100",
        1926 => x"032c8100",
        1927 => x"832c4100",
        1928 => x"032d0100",
        1929 => x"13010103",
        1930 => x"67800000",
        1931 => x"832a0b00",
        1932 => x"032d4b00",
        1933 => x"130b8b00",
        1934 => x"03298400",
        1935 => x"832c0400",
        1936 => x"e3060dfe",
        1937 => x"63642d09",
        1938 => x"8357c400",
        1939 => x"13f70748",
        1940 => x"630e0706",
        1941 => x"83244401",
        1942 => x"83250401",
        1943 => x"b3849b02",
        1944 => x"b38cbc40",
        1945 => x"13871c00",
        1946 => x"3307a701",
        1947 => x"b3c48403",
        1948 => x"63f4e400",
        1949 => x"93040700",
        1950 => x"93f70740",
        1951 => x"638c070a",
        1952 => x"93850400",
        1953 => x"13050a00",
        1954 => x"ef005049",
        1955 => x"13090500",
        1956 => x"6302050c",
        1957 => x"83250401",
        1958 => x"13860c00",
        1959 => x"eff05f97",
        1960 => x"8357c400",
        1961 => x"93f7f7b7",
        1962 => x"93e70708",
        1963 => x"2316f400",
        1964 => x"23282401",
        1965 => x"232a9400",
        1966 => x"33099901",
        1967 => x"b3849441",
        1968 => x"23202401",
        1969 => x"23249400",
        1970 => x"13090d00",
        1971 => x"63742d01",
        1972 => x"13090d00",
        1973 => x"03250400",
        1974 => x"93850a00",
        1975 => x"13060900",
        1976 => x"eff01f97",
        1977 => x"83278400",
        1978 => x"b38aaa01",
        1979 => x"b3872741",
        1980 => x"2324f400",
        1981 => x"83270400",
        1982 => x"b3872701",
        1983 => x"2320f400",
        1984 => x"83a78900",
        1985 => x"b387a741",
        1986 => x"23a4f900",
        1987 => x"e38007ee",
        1988 => x"130d0000",
        1989 => x"6ff05ff2",
        1990 => x"130a0500",
        1991 => x"13840500",
        1992 => x"930a0000",
        1993 => x"130d0000",
        1994 => x"930b3000",
        1995 => x"130c2000",
        1996 => x"6ff09ff0",
        1997 => x"13860400",
        1998 => x"13050a00",
        1999 => x"ef001053",
        2000 => x"13090500",
        2001 => x"e31605f6",
        2002 => x"83250401",
        2003 => x"13050a00",
        2004 => x"ef00502d",
        2005 => x"9307c000",
        2006 => x"2320fa00",
        2007 => x"8357c400",
        2008 => x"1305f0ff",
        2009 => x"93e70704",
        2010 => x"2316f400",
        2011 => x"23a40900",
        2012 => x"6ff01fe8",
        2013 => x"83d7c500",
        2014 => x"130101f5",
        2015 => x"2324810a",
        2016 => x"2322910a",
        2017 => x"2320210b",
        2018 => x"232c4109",
        2019 => x"2326110a",
        2020 => x"232e3109",
        2021 => x"232a5109",
        2022 => x"23286109",
        2023 => x"23267109",
        2024 => x"23248109",
        2025 => x"23229109",
        2026 => x"2320a109",
        2027 => x"232eb107",
        2028 => x"93f70708",
        2029 => x"130a0500",
        2030 => x"13890500",
        2031 => x"93040600",
        2032 => x"13840600",
        2033 => x"63880706",
        2034 => x"83a70501",
        2035 => x"63940706",
        2036 => x"93050004",
        2037 => x"ef009034",
        2038 => x"2320a900",
        2039 => x"2328a900",
        2040 => x"63160504",
        2041 => x"9307c000",
        2042 => x"2320fa00",
        2043 => x"1305f0ff",
        2044 => x"8320c10a",
        2045 => x"0324810a",
        2046 => x"8324410a",
        2047 => x"0329010a",
        2048 => x"8329c109",
        2049 => x"032a8109",
        2050 => x"832a4109",
        2051 => x"032b0109",
        2052 => x"832bc108",
        2053 => x"032c8108",
        2054 => x"832c4108",
        2055 => x"032d0108",
        2056 => x"832dc107",
        2057 => x"1301010b",
        2058 => x"67800000",
        2059 => x"93070004",
        2060 => x"232af900",
        2061 => x"93070002",
        2062 => x"a304f102",
        2063 => x"93070003",
        2064 => x"23220102",
        2065 => x"2305f102",
        2066 => x"23268100",
        2067 => x"930c5002",
        2068 => x"373b0000",
        2069 => x"b73b0000",
        2070 => x"373d0000",
        2071 => x"372c0000",
        2072 => x"930a0000",
        2073 => x"13840400",
        2074 => x"83470400",
        2075 => x"63840700",
        2076 => x"639c970d",
        2077 => x"b30d9440",
        2078 => x"63069402",
        2079 => x"93860d00",
        2080 => x"13860400",
        2081 => x"93050900",
        2082 => x"13050a00",
        2083 => x"eff09fbb",
        2084 => x"9307f0ff",
        2085 => x"6306f524",
        2086 => x"83274102",
        2087 => x"b387b701",
        2088 => x"2322f102",
        2089 => x"83470400",
        2090 => x"638c0722",
        2091 => x"9307f0ff",
        2092 => x"93041400",
        2093 => x"23280100",
        2094 => x"232e0100",
        2095 => x"232af100",
        2096 => x"232c0100",
        2097 => x"a3090104",
        2098 => x"23240106",
        2099 => x"930d1000",
        2100 => x"83c50400",
        2101 => x"13065000",
        2102 => x"13058b28",
        2103 => x"ef005012",
        2104 => x"83270101",
        2105 => x"13841400",
        2106 => x"63140506",
        2107 => x"13f70701",
        2108 => x"63060700",
        2109 => x"13070002",
        2110 => x"a309e104",
        2111 => x"13f78700",
        2112 => x"63060700",
        2113 => x"1307b002",
        2114 => x"a309e104",
        2115 => x"83c60400",
        2116 => x"1307a002",
        2117 => x"638ce604",
        2118 => x"8327c101",
        2119 => x"13840400",
        2120 => x"93060000",
        2121 => x"13069000",
        2122 => x"1305a000",
        2123 => x"03470400",
        2124 => x"93051400",
        2125 => x"130707fd",
        2126 => x"637ce608",
        2127 => x"63840604",
        2128 => x"232ef100",
        2129 => x"6f000004",
        2130 => x"13041400",
        2131 => x"6ff0dff1",
        2132 => x"13078b28",
        2133 => x"3305e540",
        2134 => x"3395ad00",
        2135 => x"b3e7a700",
        2136 => x"2328f100",
        2137 => x"93040400",
        2138 => x"6ff09ff6",
        2139 => x"0327c100",
        2140 => x"93064700",
        2141 => x"03270700",
        2142 => x"2326d100",
        2143 => x"63400704",
        2144 => x"232ee100",
        2145 => x"03470400",
        2146 => x"9307e002",
        2147 => x"6316f708",
        2148 => x"03471400",
        2149 => x"9307a002",
        2150 => x"631af704",
        2151 => x"8327c100",
        2152 => x"13042400",
        2153 => x"13874700",
        2154 => x"83a70700",
        2155 => x"2326e100",
        2156 => x"63ca0702",
        2157 => x"232af100",
        2158 => x"6f000006",
        2159 => x"3307e040",
        2160 => x"93e72700",
        2161 => x"232ee100",
        2162 => x"2328f100",
        2163 => x"6ff09ffb",
        2164 => x"b387a702",
        2165 => x"13840500",
        2166 => x"93061000",
        2167 => x"b387e700",
        2168 => x"6ff0dff4",
        2169 => x"9307f0ff",
        2170 => x"6ff0dffc",
        2171 => x"13041400",
        2172 => x"232a0100",
        2173 => x"93060000",
        2174 => x"93070000",
        2175 => x"13069000",
        2176 => x"1305a000",
        2177 => x"03470400",
        2178 => x"93051400",
        2179 => x"130707fd",
        2180 => x"6372e608",
        2181 => x"e39006fa",
        2182 => x"83450400",
        2183 => x"13063000",
        2184 => x"13850b29",
        2185 => x"ef00c07d",
        2186 => x"63020502",
        2187 => x"93870b29",
        2188 => x"3305f540",
        2189 => x"83270101",
        2190 => x"13070004",
        2191 => x"3317a700",
        2192 => x"b3e7e700",
        2193 => x"13041400",
        2194 => x"2328f100",
        2195 => x"83450400",
        2196 => x"13066000",
        2197 => x"13054d29",
        2198 => x"93041400",
        2199 => x"2304b102",
        2200 => x"ef00007a",
        2201 => x"630a0508",
        2202 => x"63980a04",
        2203 => x"03270101",
        2204 => x"8327c100",
        2205 => x"13770710",
        2206 => x"63080702",
        2207 => x"93874700",
        2208 => x"2326f100",
        2209 => x"83274102",
        2210 => x"b3873701",
        2211 => x"2322f102",
        2212 => x"6ff05fdd",
        2213 => x"b387a702",
        2214 => x"13840500",
        2215 => x"93061000",
        2216 => x"b387e700",
        2217 => x"6ff01ff6",
        2218 => x"93877700",
        2219 => x"93f787ff",
        2220 => x"93878700",
        2221 => x"6ff0dffc",
        2222 => x"1307c100",
        2223 => x"93064cc4",
        2224 => x"13060900",
        2225 => x"93050101",
        2226 => x"13050a00",
        2227 => x"97000000",
        2228 => x"e7000000",
        2229 => x"9307f0ff",
        2230 => x"93090500",
        2231 => x"e314f5fa",
        2232 => x"8357c900",
        2233 => x"1305f0ff",
        2234 => x"93f70704",
        2235 => x"e39207d0",
        2236 => x"03254102",
        2237 => x"6ff0dfcf",
        2238 => x"1307c100",
        2239 => x"93064cc4",
        2240 => x"13060900",
        2241 => x"93050101",
        2242 => x"13050a00",
        2243 => x"ef00801b",
        2244 => x"6ff05ffc",
        2245 => x"130101fd",
        2246 => x"232c4101",
        2247 => x"83a70501",
        2248 => x"130a0700",
        2249 => x"03a78500",
        2250 => x"23248102",
        2251 => x"23202103",
        2252 => x"232e3101",
        2253 => x"232a5101",
        2254 => x"23261102",
        2255 => x"23229102",
        2256 => x"23286101",
        2257 => x"23267101",
        2258 => x"93090500",
        2259 => x"13840500",
        2260 => x"13090600",
        2261 => x"938a0600",
        2262 => x"63d4e700",
        2263 => x"93070700",
        2264 => x"2320f900",
        2265 => x"03473404",
        2266 => x"63060700",
        2267 => x"93871700",
        2268 => x"2320f900",
        2269 => x"83270400",
        2270 => x"93f70702",
        2271 => x"63880700",
        2272 => x"83270900",
        2273 => x"93872700",
        2274 => x"2320f900",
        2275 => x"83240400",
        2276 => x"93f46400",
        2277 => x"639e0400",
        2278 => x"130b9401",
        2279 => x"930bf0ff",
        2280 => x"8327c400",
        2281 => x"03270900",
        2282 => x"b387e740",
        2283 => x"63c2f408",
        2284 => x"83473404",
        2285 => x"b336f000",
        2286 => x"83270400",
        2287 => x"93f70702",
        2288 => x"6390070c",
        2289 => x"13063404",
        2290 => x"93850a00",
        2291 => x"13850900",
        2292 => x"e7000a00",
        2293 => x"9307f0ff",
        2294 => x"6308f506",
        2295 => x"83270400",
        2296 => x"13074000",
        2297 => x"93040000",
        2298 => x"93f76700",
        2299 => x"639ce700",
        2300 => x"8324c400",
        2301 => x"83270900",
        2302 => x"b384f440",
        2303 => x"63d40400",
        2304 => x"93040000",
        2305 => x"83278400",
        2306 => x"03270401",
        2307 => x"6356f700",
        2308 => x"b387e740",
        2309 => x"b384f400",
        2310 => x"13090000",
        2311 => x"1304a401",
        2312 => x"130bf0ff",
        2313 => x"63902409",
        2314 => x"13050000",
        2315 => x"6f000002",
        2316 => x"93061000",
        2317 => x"13060b00",
        2318 => x"93850a00",
        2319 => x"13850900",
        2320 => x"e7000a00",
        2321 => x"631a7503",
        2322 => x"1305f0ff",
        2323 => x"8320c102",
        2324 => x"03248102",
        2325 => x"83244102",
        2326 => x"03290102",
        2327 => x"8329c101",
        2328 => x"032a8101",
        2329 => x"832a4101",
        2330 => x"032b0101",
        2331 => x"832bc100",
        2332 => x"13010103",
        2333 => x"67800000",
        2334 => x"93841400",
        2335 => x"6ff05ff2",
        2336 => x"3307d400",
        2337 => x"13060003",
        2338 => x"a301c704",
        2339 => x"03475404",
        2340 => x"93871600",
        2341 => x"b307f400",
        2342 => x"93862600",
        2343 => x"a381e704",
        2344 => x"6ff05ff2",
        2345 => x"93061000",
        2346 => x"13060400",
        2347 => x"93850a00",
        2348 => x"13850900",
        2349 => x"e7000a00",
        2350 => x"e30865f9",
        2351 => x"13091900",
        2352 => x"6ff05ff6",
        2353 => x"130101fd",
        2354 => x"23248102",
        2355 => x"23229102",
        2356 => x"23202103",
        2357 => x"232e3101",
        2358 => x"23261102",
        2359 => x"232c4101",
        2360 => x"232a5101",
        2361 => x"23286101",
        2362 => x"83c88501",
        2363 => x"93078007",
        2364 => x"93040500",
        2365 => x"13840500",
        2366 => x"13090600",
        2367 => x"93890600",
        2368 => x"63ee1701",
        2369 => x"93072006",
        2370 => x"93863504",
        2371 => x"63ee1701",
        2372 => x"63840828",
        2373 => x"93078005",
        2374 => x"6388f822",
        2375 => x"930a2404",
        2376 => x"23011405",
        2377 => x"6f004004",
        2378 => x"9387d8f9",
        2379 => x"93f7f70f",
        2380 => x"13065001",
        2381 => x"e364f6fe",
        2382 => x"37360000",
        2383 => x"93972700",
        2384 => x"1306462c",
        2385 => x"b387c700",
        2386 => x"83a70700",
        2387 => x"67800700",
        2388 => x"83270700",
        2389 => x"938a2504",
        2390 => x"93864700",
        2391 => x"83a70700",
        2392 => x"2320d700",
        2393 => x"2381f504",
        2394 => x"93071000",
        2395 => x"6f008026",
        2396 => x"83a70500",
        2397 => x"03250700",
        2398 => x"13f60708",
        2399 => x"93054500",
        2400 => x"63060602",
        2401 => x"83270500",
        2402 => x"2320b700",
        2403 => x"37380000",
        2404 => x"63d80700",
        2405 => x"1307d002",
        2406 => x"b307f040",
        2407 => x"a301e404",
        2408 => x"1308c829",
        2409 => x"1307a000",
        2410 => x"6f008006",
        2411 => x"13f60704",
        2412 => x"83270500",
        2413 => x"2320b700",
        2414 => x"e30a06fc",
        2415 => x"93970701",
        2416 => x"93d70741",
        2417 => x"6ff09ffc",
        2418 => x"03a60500",
        2419 => x"83270700",
        2420 => x"13750608",
        2421 => x"93854700",
        2422 => x"63080500",
        2423 => x"2320b700",
        2424 => x"83a70700",
        2425 => x"6f004001",
        2426 => x"13760604",
        2427 => x"2320b700",
        2428 => x"e30806fe",
        2429 => x"83d70700",
        2430 => x"37380000",
        2431 => x"1307f006",
        2432 => x"1308c829",
        2433 => x"6388e814",
        2434 => x"1307a000",
        2435 => x"a3010404",
        2436 => x"03264400",
        2437 => x"2324c400",
        2438 => x"63480600",
        2439 => x"83250400",
        2440 => x"93f5b5ff",
        2441 => x"2320b400",
        2442 => x"63960700",
        2443 => x"938a0600",
        2444 => x"63040602",
        2445 => x"938a0600",
        2446 => x"33f6e702",
        2447 => x"938afaff",
        2448 => x"3306c800",
        2449 => x"03460600",
        2450 => x"2380ca00",
        2451 => x"13860700",
        2452 => x"b3d7e702",
        2453 => x"e372e6fe",
        2454 => x"93078000",
        2455 => x"6314f702",
        2456 => x"83270400",
        2457 => x"93f71700",
        2458 => x"638e0700",
        2459 => x"03274400",
        2460 => x"83270401",
        2461 => x"63c8e700",
        2462 => x"93070003",
        2463 => x"a38ffafe",
        2464 => x"938afaff",
        2465 => x"b3865641",
        2466 => x"2328d400",
        2467 => x"13870900",
        2468 => x"93060900",
        2469 => x"1306c100",
        2470 => x"93050400",
        2471 => x"13850400",
        2472 => x"eff05fc7",
        2473 => x"130af0ff",
        2474 => x"631c4513",
        2475 => x"1305f0ff",
        2476 => x"8320c102",
        2477 => x"03248102",
        2478 => x"83244102",
        2479 => x"03290102",
        2480 => x"8329c101",
        2481 => x"032a8101",
        2482 => x"832a4101",
        2483 => x"032b0101",
        2484 => x"13010103",
        2485 => x"67800000",
        2486 => x"83a70500",
        2487 => x"93e70702",
        2488 => x"23a0f500",
        2489 => x"37380000",
        2490 => x"93088007",
        2491 => x"1308082b",
        2492 => x"a3021405",
        2493 => x"03260400",
        2494 => x"83250700",
        2495 => x"13750608",
        2496 => x"83a70500",
        2497 => x"93854500",
        2498 => x"631a0500",
        2499 => x"13750604",
        2500 => x"63060500",
        2501 => x"93970701",
        2502 => x"93d70701",
        2503 => x"2320b700",
        2504 => x"13771600",
        2505 => x"63060700",
        2506 => x"13660602",
        2507 => x"2320c400",
        2508 => x"13070001",
        2509 => x"e39c07ec",
        2510 => x"03260400",
        2511 => x"1376f6fd",
        2512 => x"2320c400",
        2513 => x"6ff09fec",
        2514 => x"37380000",
        2515 => x"1308c829",
        2516 => x"6ff01ffa",
        2517 => x"13078000",
        2518 => x"6ff05feb",
        2519 => x"03a60500",
        2520 => x"83270700",
        2521 => x"83a54501",
        2522 => x"13780608",
        2523 => x"13854700",
        2524 => x"630a0800",
        2525 => x"2320a700",
        2526 => x"83a70700",
        2527 => x"23a0b700",
        2528 => x"6f008001",
        2529 => x"2320a700",
        2530 => x"13760604",
        2531 => x"83a70700",
        2532 => x"e30606fe",
        2533 => x"2390b700",
        2534 => x"23280400",
        2535 => x"938a0600",
        2536 => x"6ff0dfee",
        2537 => x"83270700",
        2538 => x"03a64500",
        2539 => x"93050000",
        2540 => x"93864700",
        2541 => x"2320d700",
        2542 => x"83aa0700",
        2543 => x"13850a00",
        2544 => x"ef000024",
        2545 => x"63060500",
        2546 => x"33055541",
        2547 => x"2322a400",
        2548 => x"83274400",
        2549 => x"2328f400",
        2550 => x"a3010404",
        2551 => x"6ff01feb",
        2552 => x"83260401",
        2553 => x"13860a00",
        2554 => x"93050900",
        2555 => x"13850400",
        2556 => x"e7800900",
        2557 => x"e30c45eb",
        2558 => x"83270400",
        2559 => x"93f72700",
        2560 => x"63940704",
        2561 => x"8327c100",
        2562 => x"0325c400",
        2563 => x"e352f5ea",
        2564 => x"13850700",
        2565 => x"6ff0dfe9",
        2566 => x"93061000",
        2567 => x"13860a00",
        2568 => x"93050900",
        2569 => x"13850400",
        2570 => x"e7800900",
        2571 => x"e30065e9",
        2572 => x"130a1a00",
        2573 => x"8327c400",
        2574 => x"0327c100",
        2575 => x"b387e740",
        2576 => x"e34cfafc",
        2577 => x"6ff01ffc",
        2578 => x"130a0000",
        2579 => x"930a9401",
        2580 => x"130bf0ff",
        2581 => x"6ff01ffe",
        2582 => x"130101ff",
        2583 => x"23248100",
        2584 => x"13840500",
        2585 => x"83a50500",
        2586 => x"23229100",
        2587 => x"23261100",
        2588 => x"93040500",
        2589 => x"63840500",
        2590 => x"eff01ffe",
        2591 => x"93050400",
        2592 => x"03248100",
        2593 => x"8320c100",
        2594 => x"13850400",
        2595 => x"83244100",
        2596 => x"13010101",
        2597 => x"6f000019",
        2598 => x"83a7c187",
        2599 => x"6380a716",
        2600 => x"83274502",
        2601 => x"130101fe",
        2602 => x"232c8100",
        2603 => x"232e1100",
        2604 => x"232a9100",
        2605 => x"23282101",
        2606 => x"23263101",
        2607 => x"13040500",
        2608 => x"63840702",
        2609 => x"83a7c700",
        2610 => x"93040000",
        2611 => x"13090008",
        2612 => x"6392070e",
        2613 => x"83274402",
        2614 => x"83a50700",
        2615 => x"63860500",
        2616 => x"13050400",
        2617 => x"ef000014",
        2618 => x"83254401",
        2619 => x"63860500",
        2620 => x"13050400",
        2621 => x"ef000013",
        2622 => x"83254402",
        2623 => x"63860500",
        2624 => x"13050400",
        2625 => x"ef000012",
        2626 => x"83258403",
        2627 => x"63860500",
        2628 => x"13050400",
        2629 => x"ef000011",
        2630 => x"8325c403",
        2631 => x"63860500",
        2632 => x"13050400",
        2633 => x"ef000010",
        2634 => x"83250404",
        2635 => x"63860500",
        2636 => x"13050400",
        2637 => x"ef00000f",
        2638 => x"8325c405",
        2639 => x"63860500",
        2640 => x"13050400",
        2641 => x"ef00000e",
        2642 => x"83258405",
        2643 => x"63860500",
        2644 => x"13050400",
        2645 => x"ef00000d",
        2646 => x"83254403",
        2647 => x"63860500",
        2648 => x"13050400",
        2649 => x"ef00000c",
        2650 => x"83278401",
        2651 => x"638a0706",
        2652 => x"83278402",
        2653 => x"13050400",
        2654 => x"e7800700",
        2655 => x"83258404",
        2656 => x"63800506",
        2657 => x"13050400",
        2658 => x"03248101",
        2659 => x"8320c101",
        2660 => x"83244101",
        2661 => x"03290101",
        2662 => x"8329c100",
        2663 => x"13010102",
        2664 => x"6ff09feb",
        2665 => x"b3859500",
        2666 => x"83a50500",
        2667 => x"63900502",
        2668 => x"93844400",
        2669 => x"83274402",
        2670 => x"83a5c700",
        2671 => x"e39424ff",
        2672 => x"13050400",
        2673 => x"ef000006",
        2674 => x"6ff0dff0",
        2675 => x"83a90500",
        2676 => x"13050400",
        2677 => x"ef000005",
        2678 => x"93850900",
        2679 => x"6ff01ffd",
        2680 => x"8320c101",
        2681 => x"03248101",
        2682 => x"83244101",
        2683 => x"03290101",
        2684 => x"8329c100",
        2685 => x"13010102",
        2686 => x"67800000",
        2687 => x"67800000",
        2688 => x"93f5f50f",
        2689 => x"3306c500",
        2690 => x"6316c500",
        2691 => x"13050000",
        2692 => x"67800000",
        2693 => x"83470500",
        2694 => x"e38cb7fe",
        2695 => x"13051500",
        2696 => x"6ff09ffe",
        2697 => x"638a050e",
        2698 => x"83a7c5ff",
        2699 => x"130101fe",
        2700 => x"232c8100",
        2701 => x"232e1100",
        2702 => x"1384c5ff",
        2703 => x"63d40700",
        2704 => x"3304f400",
        2705 => x"2326a100",
        2706 => x"ef000034",
        2707 => x"83a78188",
        2708 => x"0325c100",
        2709 => x"639e0700",
        2710 => x"23220400",
        2711 => x"23a48188",
        2712 => x"03248101",
        2713 => x"8320c101",
        2714 => x"13010102",
        2715 => x"6f000032",
        2716 => x"6374f402",
        2717 => x"03260400",
        2718 => x"b306c400",
        2719 => x"639ad700",
        2720 => x"83a60700",
        2721 => x"83a74700",
        2722 => x"b386c600",
        2723 => x"2320d400",
        2724 => x"2322f400",
        2725 => x"6ff09ffc",
        2726 => x"13870700",
        2727 => x"83a74700",
        2728 => x"63840700",
        2729 => x"e37af4fe",
        2730 => x"83260700",
        2731 => x"3306d700",
        2732 => x"63188602",
        2733 => x"03260400",
        2734 => x"b386c600",
        2735 => x"2320d700",
        2736 => x"3306d700",
        2737 => x"e39ec7f8",
        2738 => x"03a60700",
        2739 => x"83a74700",
        2740 => x"b306d600",
        2741 => x"2320d700",
        2742 => x"2322f700",
        2743 => x"6ff05ff8",
        2744 => x"6378c400",
        2745 => x"9307c000",
        2746 => x"2320f500",
        2747 => x"6ff05ff7",
        2748 => x"03260400",
        2749 => x"b306c400",
        2750 => x"639ad700",
        2751 => x"83a60700",
        2752 => x"83a74700",
        2753 => x"b386c600",
        2754 => x"2320d400",
        2755 => x"2322f400",
        2756 => x"23228700",
        2757 => x"6ff0dff4",
        2758 => x"67800000",
        2759 => x"130101fe",
        2760 => x"232a9100",
        2761 => x"93843500",
        2762 => x"93f4c4ff",
        2763 => x"23282101",
        2764 => x"232e1100",
        2765 => x"232c8100",
        2766 => x"23263101",
        2767 => x"93848400",
        2768 => x"9307c000",
        2769 => x"13090500",
        2770 => x"63f4f406",
        2771 => x"9304c000",
        2772 => x"63e2b406",
        2773 => x"13050900",
        2774 => x"ef000023",
        2775 => x"03a78188",
        2776 => x"93868188",
        2777 => x"13040700",
        2778 => x"631a0406",
        2779 => x"1384c188",
        2780 => x"83270400",
        2781 => x"639a0700",
        2782 => x"93050000",
        2783 => x"13050900",
        2784 => x"ef00001c",
        2785 => x"2320a400",
        2786 => x"93850400",
        2787 => x"13050900",
        2788 => x"ef00001b",
        2789 => x"9309f0ff",
        2790 => x"631a350b",
        2791 => x"9307c000",
        2792 => x"2320f900",
        2793 => x"13050900",
        2794 => x"ef00401e",
        2795 => x"6f000001",
        2796 => x"e3d004fa",
        2797 => x"9307c000",
        2798 => x"2320f900",
        2799 => x"13050000",
        2800 => x"8320c101",
        2801 => x"03248101",
        2802 => x"83244101",
        2803 => x"03290101",
        2804 => x"8329c100",
        2805 => x"13010102",
        2806 => x"67800000",
        2807 => x"83270400",
        2808 => x"b3879740",
        2809 => x"63ce0704",
        2810 => x"1306b000",
        2811 => x"637af600",
        2812 => x"2320f400",
        2813 => x"3304f400",
        2814 => x"23209400",
        2815 => x"6f000001",
        2816 => x"83274400",
        2817 => x"631a8702",
        2818 => x"23a0f600",
        2819 => x"13050900",
        2820 => x"ef00c017",
        2821 => x"1305b400",
        2822 => x"93074400",
        2823 => x"137585ff",
        2824 => x"3307f540",
        2825 => x"e30ef5f8",
        2826 => x"3304e400",
        2827 => x"b387a740",
        2828 => x"2320f400",
        2829 => x"6ff0dff8",
        2830 => x"2322f700",
        2831 => x"6ff01ffd",
        2832 => x"13070400",
        2833 => x"03244400",
        2834 => x"6ff01ff2",
        2835 => x"13043500",
        2836 => x"1374c4ff",
        2837 => x"e30285fa",
        2838 => x"b305a440",
        2839 => x"13050900",
        2840 => x"ef00000e",
        2841 => x"e31a35f9",
        2842 => x"6ff05ff3",
        2843 => x"130101fe",
        2844 => x"232c8100",
        2845 => x"232e1100",
        2846 => x"232a9100",
        2847 => x"23282101",
        2848 => x"23263101",
        2849 => x"23244101",
        2850 => x"13040600",
        2851 => x"63940502",
        2852 => x"03248101",
        2853 => x"8320c101",
        2854 => x"83244101",
        2855 => x"03290101",
        2856 => x"8329c100",
        2857 => x"032a8100",
        2858 => x"93050600",
        2859 => x"13010102",
        2860 => x"6ff0dfe6",
        2861 => x"63180602",
        2862 => x"eff0dfd6",
        2863 => x"93040000",
        2864 => x"8320c101",
        2865 => x"03248101",
        2866 => x"03290101",
        2867 => x"8329c100",
        2868 => x"032a8100",
        2869 => x"13850400",
        2870 => x"83244101",
        2871 => x"13010102",
        2872 => x"67800000",
        2873 => x"130a0500",
        2874 => x"13890500",
        2875 => x"ef00400a",
        2876 => x"93090500",
        2877 => x"63688500",
        2878 => x"93571500",
        2879 => x"93040900",
        2880 => x"e3e087fc",
        2881 => x"93050400",
        2882 => x"13050a00",
        2883 => x"eff01fe1",
        2884 => x"93040500",
        2885 => x"e30605fa",
        2886 => x"13060400",
        2887 => x"63f48900",
        2888 => x"13860900",
        2889 => x"93050900",
        2890 => x"13850400",
        2891 => x"efe05fae",
        2892 => x"93050900",
        2893 => x"13050a00",
        2894 => x"eff0dfce",
        2895 => x"6ff05ff8",
        2896 => x"130101ff",
        2897 => x"23248100",
        2898 => x"23229100",
        2899 => x"13040500",
        2900 => x"13850500",
        2901 => x"23261100",
        2902 => x"23a20188",
        2903 => x"ef00000c",
        2904 => x"9307f0ff",
        2905 => x"6318f500",
        2906 => x"83a74188",
        2907 => x"63840700",
        2908 => x"2320f400",
        2909 => x"8320c100",
        2910 => x"03248100",
        2911 => x"83244100",
        2912 => x"13010101",
        2913 => x"67800000",
        2914 => x"67800000",
        2915 => x"67800000",
        2916 => x"83a7c5ff",
        2917 => x"1385c7ff",
        2918 => x"63d80700",
        2919 => x"b385a500",
        2920 => x"83a70500",
        2921 => x"3305f500",
        2922 => x"67800000",
        2923 => x"9308d005",
        2924 => x"73000000",
        2925 => x"63520502",
        2926 => x"130101ff",
        2927 => x"23248100",
        2928 => x"13040500",
        2929 => x"23261100",
        2930 => x"33048040",
        2931 => x"efe05fc6",
        2932 => x"23208500",
        2933 => x"6f000000",
        2934 => x"6f000000",
        2935 => x"130101ff",
        2936 => x"23261100",
        2937 => x"23248100",
        2938 => x"9308900a",
        2939 => x"73000000",
        2940 => x"13040500",
        2941 => x"635a0500",
        2942 => x"33048040",
        2943 => x"efe05fc3",
        2944 => x"23208500",
        2945 => x"1304f0ff",
        2946 => x"8320c100",
        2947 => x"13050400",
        2948 => x"03248100",
        2949 => x"13010101",
        2950 => x"67800000",
        2951 => x"83a70189",
        2952 => x"130101ff",
        2953 => x"23261100",
        2954 => x"93060500",
        2955 => x"13870189",
        2956 => x"639c0702",
        2957 => x"9308600d",
        2958 => x"13050000",
        2959 => x"73000000",
        2960 => x"9307f0ff",
        2961 => x"6310f502",
        2962 => x"efe09fbe",
        2963 => x"9307c000",
        2964 => x"2320f500",
        2965 => x"1305f0ff",
        2966 => x"8320c100",
        2967 => x"13010101",
        2968 => x"67800000",
        2969 => x"2320a700",
        2970 => x"83270700",
        2971 => x"9308600d",
        2972 => x"b386f600",
        2973 => x"13850600",
        2974 => x"73000000",
        2975 => x"e316d5fc",
        2976 => x"2320a700",
        2977 => x"13850700",
        2978 => x"6ff01ffd",
        2979 => x"10000000",
        2980 => x"00000000",
        2981 => x"037a5200",
        2982 => x"017c0101",
        2983 => x"1b0d0200",
        2984 => x"10000000",
        2985 => x"18000000",
        2986 => x"8cd8ffff",
        2987 => x"78040000",
        2988 => x"00000000",
        2989 => x"10000000",
        2990 => x"00000000",
        2991 => x"037a5200",
        2992 => x"017c0101",
        2993 => x"1b0d0200",
        2994 => x"10000000",
        2995 => x"18000000",
        2996 => x"dcdcffff",
        2997 => x"50040000",
        2998 => x"00000000",
        2999 => x"10000000",
        3000 => x"00000000",
        3001 => x"037a5200",
        3002 => x"017c0101",
        3003 => x"1b0d0200",
        3004 => x"10000000",
        3005 => x"18000000",
        3006 => x"04e1ffff",
        3007 => x"30040000",
        3008 => x"00000000",
        3009 => x"10000000",
        3010 => x"00000000",
        3011 => x"037a5200",
        3012 => x"017c0101",
        3013 => x"1b0d0200",
        3014 => x"10000000",
        3015 => x"18000000",
        3016 => x"0ce5ffff",
        3017 => x"e4030000",
        3018 => x"00000000",
        3019 => x"2c020000",
        3020 => x"9c010000",
        3021 => x"9c010000",
        3022 => x"9c010000",
        3023 => x"9c010000",
        3024 => x"10020000",
        3025 => x"9c010000",
        3026 => x"d0010000",
        3027 => x"9c010000",
        3028 => x"9c010000",
        3029 => x"d0010000",
        3030 => x"9c010000",
        3031 => x"9c010000",
        3032 => x"9c010000",
        3033 => x"9c010000",
        3034 => x"9c010000",
        3035 => x"9c010000",
        3036 => x"9c010000",
        3037 => x"80010000",
        3038 => x"28040000",
        3039 => x"28040000",
        3040 => x"28040000",
        3041 => x"80040000",
        3042 => x"28040000",
        3043 => x"28040000",
        3044 => x"28040000",
        3045 => x"28040000",
        3046 => x"28040000",
        3047 => x"28040000",
        3048 => x"28040000",
        3049 => x"48040000",
        3050 => x"ec040000",
        3051 => x"b4040000",
        3052 => x"b4040000",
        3053 => x"b4040000",
        3054 => x"b4040000",
        3055 => x"e0040000",
        3056 => x"74050000",
        3057 => x"4c050000",
        3058 => x"b4040000",
        3059 => x"b4040000",
        3060 => x"b4040000",
        3061 => x"b4040000",
        3062 => x"b4040000",
        3063 => x"b4040000",
        3064 => x"b4040000",
        3065 => x"b4040000",
        3066 => x"b4040000",
        3067 => x"b4040000",
        3068 => x"b4040000",
        3069 => x"b4040000",
        3070 => x"b4040000",
        3071 => x"b4040000",
        3072 => x"cc040000",
        3073 => x"cc040000",
        3074 => x"b4040000",
        3075 => x"b4040000",
        3076 => x"b4040000",
        3077 => x"b4040000",
        3078 => x"b4040000",
        3079 => x"b4040000",
        3080 => x"b4040000",
        3081 => x"b4040000",
        3082 => x"b4040000",
        3083 => x"b4040000",
        3084 => x"b4040000",
        3085 => x"b4040000",
        3086 => x"e0040000",
        3087 => x"ec040000",
        3088 => x"04050000",
        3089 => x"34050000",
        3090 => x"b4040000",
        3091 => x"b4040000",
        3092 => x"b4040000",
        3093 => x"b4040000",
        3094 => x"b4040000",
        3095 => x"b4040000",
        3096 => x"1c050000",
        3097 => x"b4040000",
        3098 => x"b4040000",
        3099 => x"b4040000",
        3100 => x"b4040000",
        3101 => x"cc040000",
        3102 => x"cc040000",
        3103 => x"00010202",
        3104 => x"03030303",
        3105 => x"04040404",
        3106 => x"04040404",
        3107 => x"05050505",
        3108 => x"05050505",
        3109 => x"05050505",
        3110 => x"05050505",
        3111 => x"06060606",
        3112 => x"06060606",
        3113 => x"06060606",
        3114 => x"06060606",
        3115 => x"06060606",
        3116 => x"06060606",
        3117 => x"06060606",
        3118 => x"06060606",
        3119 => x"07070707",
        3120 => x"07070707",
        3121 => x"07070707",
        3122 => x"07070707",
        3123 => x"07070707",
        3124 => x"07070707",
        3125 => x"07070707",
        3126 => x"07070707",
        3127 => x"07070707",
        3128 => x"07070707",
        3129 => x"07070707",
        3130 => x"07070707",
        3131 => x"07070707",
        3132 => x"07070707",
        3133 => x"07070707",
        3134 => x"07070707",
        3135 => x"08080808",
        3136 => x"08080808",
        3137 => x"08080808",
        3138 => x"08080808",
        3139 => x"08080808",
        3140 => x"08080808",
        3141 => x"08080808",
        3142 => x"08080808",
        3143 => x"08080808",
        3144 => x"08080808",
        3145 => x"08080808",
        3146 => x"08080808",
        3147 => x"08080808",
        3148 => x"08080808",
        3149 => x"08080808",
        3150 => x"08080808",
        3151 => x"08080808",
        3152 => x"08080808",
        3153 => x"08080808",
        3154 => x"08080808",
        3155 => x"08080808",
        3156 => x"08080808",
        3157 => x"08080808",
        3158 => x"08080808",
        3159 => x"08080808",
        3160 => x"08080808",
        3161 => x"08080808",
        3162 => x"08080808",
        3163 => x"08080808",
        3164 => x"08080808",
        3165 => x"08080808",
        3166 => x"08080808",
        3167 => x"0d0a0d0a",
        3168 => x"44697370",
        3169 => x"6c617969",
        3170 => x"6e672074",
        3171 => x"68652074",
        3172 => x"696d6520",
        3173 => x"70617373",
        3174 => x"65642073",
        3175 => x"696e6365",
        3176 => x"20726573",
        3177 => x"65740d0a",
        3178 => x"0d0a0000",
        3179 => x"2530356c",
        3180 => x"643a2530",
        3181 => x"366c6420",
        3182 => x"20202530",
        3183 => x"326c643a",
        3184 => x"2530326c",
        3185 => x"643a2530",
        3186 => x"326c640d",
        3187 => x"00000000",
        3188 => x"696e7465",
        3189 => x"72727570",
        3190 => x"74000000",
        3191 => x"52495343",
        3192 => x"2d562052",
        3193 => x"56333249",
        3194 => x"4d206261",
        3195 => x"7265206d",
        3196 => x"6574616c",
        3197 => x"2070726f",
        3198 => x"63657373",
        3199 => x"6f720000",
        3200 => x"54686520",
        3201 => x"48616775",
        3202 => x"6520556e",
        3203 => x"69766572",
        3204 => x"73697479",
        3205 => x"206f6620",
        3206 => x"4170706c",
        3207 => x"69656420",
        3208 => x"53636965",
        3209 => x"6e636573",
        3210 => x"00000000",
        3211 => x"44657061",
        3212 => x"72746d65",
        3213 => x"6e74206f",
        3214 => x"6620456c",
        3215 => x"65637472",
        3216 => x"6963616c",
        3217 => x"20456e67",
        3218 => x"696e6565",
        3219 => x"72696e67",
        3220 => x"00000000",
        3221 => x"4a2e452e",
        3222 => x"4a2e206f",
        3223 => x"70206465",
        3224 => x"6e204272",
        3225 => x"6f757700",
        3226 => x"3c627265",
        3227 => x"616b3e0d",
        3228 => x"0a000000",
        3229 => x"0d0a4542",
        3230 => x"5245414b",
        3231 => x"21206d69",
        3232 => x"70203d20",
        3233 => x"00000000",
        3234 => x"232d302b",
        3235 => x"20000000",
        3236 => x"686c4c00",
        3237 => x"65666745",
        3238 => x"46470000",
        3239 => x"30313233",
        3240 => x"34353637",
        3241 => x"38394142",
        3242 => x"43444546",
        3243 => x"00000000",
        3244 => x"30313233",
        3245 => x"34353637",
        3246 => x"38396162",
        3247 => x"63646566",
        3248 => x"00000000",
        3249 => x"50250000",
        3250 => x"70250000",
        3251 => x"1c250000",
        3252 => x"1c250000",
        3253 => x"1c250000",
        3254 => x"1c250000",
        3255 => x"70250000",
        3256 => x"1c250000",
        3257 => x"1c250000",
        3258 => x"1c250000",
        3259 => x"1c250000",
        3260 => x"5c270000",
        3261 => x"c8250000",
        3262 => x"d8260000",
        3263 => x"1c250000",
        3264 => x"1c250000",
        3265 => x"a4270000",
        3266 => x"1c250000",
        3267 => x"c8250000",
        3268 => x"1c250000",
        3269 => x"1c250000",
        3270 => x"e4260000",
        3271 => x"18000020",
        3272 => x"d0310000",
        3273 => x"dc310000",
        3274 => x"00320000",
        3275 => x"2c320000",
        3276 => x"54320000",
        3277 => x"00000000",
        3278 => x"00000000",
        3279 => x"00000000",
        3280 => x"00000000",
        3281 => x"00000000",
        3282 => x"00000000",
        3283 => x"00000000",
        3284 => x"00000000",
        3285 => x"00000000",
        3286 => x"00000000",
        3287 => x"00000000",
        3288 => x"00000000",
        3289 => x"00000000",
        3290 => x"00000000",
        3291 => x"00000000",
        3292 => x"00000000",
        3293 => x"00000000",
        3294 => x"00000000",
        3295 => x"00000000",
        3296 => x"00000000",
        3297 => x"00000000",
        3298 => x"00000000",
        3299 => x"00000000",
        3300 => x"00000000",
        3301 => x"00000000",
        3302 => x"80000020",
        3303 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
