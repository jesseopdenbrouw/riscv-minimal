-- srec2vhdl table generator
-- for input file clock.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"93804186",
           5 => x"93844187",
           6 => x"b7370000",
           7 => x"1389c731",
           8 => x"6f004001",
           9 => x"23a00000",
          10 => x"93870000",
          11 => x"93804700",
          12 => x"83a70700",
          13 => x"e3e890fe",
          14 => x"b7070020",
          15 => x"93800700",
          16 => x"93844186",
          17 => x"6f004001",
          18 => x"83270900",
          19 => x"23a0f000",
          20 => x"93804000",
          21 => x"13094900",
          22 => x"e3e890fe",
          23 => x"ef105033",
          24 => x"ef00800e",
          25 => x"13050000",
          26 => x"ef10902e",
          27 => x"130101ff",
          28 => x"23268100",
          29 => x"13040101",
          30 => x"b70700f0",
          31 => x"93870702",
          32 => x"37170000",
          33 => x"13077745",
          34 => x"23a2e700",
          35 => x"13000000",
          36 => x"0324c100",
          37 => x"13010101",
          38 => x"67800000",
          39 => x"130101fe",
          40 => x"232e8100",
          41 => x"13040102",
          42 => x"2326a4fe",
          43 => x"8327c4fe",
          44 => x"13f7f70f",
          45 => x"b70700f0",
          46 => x"93870702",
          47 => x"23a0e700",
          48 => x"13000000",
          49 => x"b70700f0",
          50 => x"93870702",
          51 => x"83a7c700",
          52 => x"93f70701",
          53 => x"e38807fe",
          54 => x"13000000",
          55 => x"13000000",
          56 => x"0324c101",
          57 => x"13010102",
          58 => x"67800000",
          59 => x"130101fe",
          60 => x"232e1100",
          61 => x"232c8100",
          62 => x"13040102",
          63 => x"2326a4fe",
          64 => x"8327c4fe",
          65 => x"63880702",
          66 => x"6f00c001",
          67 => x"8327c4fe",
          68 => x"13871700",
          69 => x"2326e4fe",
          70 => x"83c70700",
          71 => x"13850700",
          72 => x"eff0dff7",
          73 => x"8327c4fe",
          74 => x"83c70700",
          75 => x"e39007fe",
          76 => x"6f008000",
          77 => x"13000000",
          78 => x"8320c101",
          79 => x"03248101",
          80 => x"13010102",
          81 => x"67800000",
          82 => x"130101f6",
          83 => x"232e1108",
          84 => x"232c8108",
          85 => x"1304010a",
          86 => x"232204f6",
          87 => x"930784f6",
          88 => x"13070006",
          89 => x"13060700",
          90 => x"93050000",
          91 => x"13850700",
          92 => x"ef10d015",
          93 => x"eff09fef",
          94 => x"b7370000",
          95 => x"13858713",
          96 => x"eff0dff6",
          97 => x"930784fc",
          98 => x"93050000",
          99 => x"13850700",
         100 => x"ef105040",
         101 => x"032784fc",
         102 => x"8327c4fc",
         103 => x"1306c003",
         104 => x"93060000",
         105 => x"13050700",
         106 => x"93850700",
         107 => x"ef00100a",
         108 => x"13070500",
         109 => x"93870500",
         110 => x"2324e4fe",
         111 => x"2326f4fe",
         112 => x"032784fc",
         113 => x"8327c4fc",
         114 => x"1306c003",
         115 => x"93060000",
         116 => x"13050700",
         117 => x"93850700",
         118 => x"ef004026",
         119 => x"13070500",
         120 => x"93870500",
         121 => x"1306c003",
         122 => x"93060000",
         123 => x"13050700",
         124 => x"93850700",
         125 => x"ef009005",
         126 => x"13070500",
         127 => x"93870500",
         128 => x"2320e4fe",
         129 => x"2322f4fe",
         130 => x"032784fc",
         131 => x"8327c4fc",
         132 => x"37160000",
         133 => x"130606e1",
         134 => x"93060000",
         135 => x"13050700",
         136 => x"93850700",
         137 => x"ef008021",
         138 => x"13070500",
         139 => x"93870500",
         140 => x"232ce4fc",
         141 => x"232ef4fc",
         142 => x"032784fc",
         143 => x"8327c4fc",
         144 => x"93050700",
         145 => x"032704fd",
         146 => x"832784fd",
         147 => x"832604fe",
         148 => x"032684fe",
         149 => x"130544f6",
         150 => x"93080600",
         151 => x"13880600",
         152 => x"93860500",
         153 => x"37360000",
         154 => x"13068615",
         155 => x"93054006",
         156 => x"ef101027",
         157 => x"930744f6",
         158 => x"13850700",
         159 => x"eff01fe7",
         160 => x"6ff05ff0",
         161 => x"130101fb",
         162 => x"23261104",
         163 => x"23248104",
         164 => x"13040105",
         165 => x"232ea4fa",
         166 => x"232cb4fa",
         167 => x"232604fe",
         168 => x"8325c4fe",
         169 => x"2324b4fe",
         170 => x"832584fe",
         171 => x"2322b4fe",
         172 => x"032844fe",
         173 => x"032584fe",
         174 => x"8325c4fe",
         175 => x"732810c8",
         176 => x"732510c0",
         177 => x"f32510c8",
         178 => x"e31ab8fe",
         179 => x"232204ff",
         180 => x"2324a4fe",
         181 => x"2326b4fe",
         182 => x"832544fe",
         183 => x"13830500",
         184 => x"93030000",
         185 => x"93170300",
         186 => x"13070000",
         187 => x"832584fe",
         188 => x"13860500",
         189 => x"93060000",
         190 => x"b365c700",
         191 => x"232cb4fc",
         192 => x"b3e7d700",
         193 => x"232ef4fc",
         194 => x"032784fd",
         195 => x"8327c4fd",
         196 => x"37460f00",
         197 => x"13060624",
         198 => x"93060000",
         199 => x"13050700",
         200 => x"93850700",
         201 => x"ef100020",
         202 => x"13070500",
         203 => x"93870500",
         204 => x"2328e4fc",
         205 => x"232af4fc",
         206 => x"032784fd",
         207 => x"8327c4fd",
         208 => x"37460f00",
         209 => x"13060624",
         210 => x"93060000",
         211 => x"13050700",
         212 => x"93850700",
         213 => x"ef001041",
         214 => x"13070500",
         215 => x"93870500",
         216 => x"2324e4fc",
         217 => x"2326f4fc",
         218 => x"032704fd",
         219 => x"8327c4fb",
         220 => x"23a4e700",
         221 => x"032784fc",
         222 => x"8327c4fc",
         223 => x"8326c4fb",
         224 => x"23a0e600",
         225 => x"23a2f600",
         226 => x"93070000",
         227 => x"13850700",
         228 => x"8320c104",
         229 => x"03248104",
         230 => x"13010105",
         231 => x"67800000",
         232 => x"130101fd",
         233 => x"23261102",
         234 => x"23248102",
         235 => x"13040103",
         236 => x"232ea4fc",
         237 => x"b7870020",
         238 => x"13870700",
         239 => x"93070040",
         240 => x"b307f740",
         241 => x"2326f4fe",
         242 => x"8327c4fe",
         243 => x"2324f4fe",
         244 => x"83a70187",
         245 => x"63960700",
         246 => x"13878187",
         247 => x"23a8e186",
         248 => x"03a70187",
         249 => x"8327c4fd",
         250 => x"b307f700",
         251 => x"032784fe",
         252 => x"637ef700",
         253 => x"ef104075",
         254 => x"13070500",
         255 => x"9307c000",
         256 => x"2320f700",
         257 => x"9307f0ff",
         258 => x"6f000002",
         259 => x"83a70187",
         260 => x"2322f4fe",
         261 => x"03a70187",
         262 => x"8327c4fd",
         263 => x"3307f700",
         264 => x"23a8e186",
         265 => x"832744fe",
         266 => x"13850700",
         267 => x"8320c102",
         268 => x"03248102",
         269 => x"13010103",
         270 => x"67800000",
         271 => x"130101fd",
         272 => x"23229102",
         273 => x"232c4101",
         274 => x"23261102",
         275 => x"23248102",
         276 => x"23202103",
         277 => x"232e3101",
         278 => x"232a5101",
         279 => x"23286101",
         280 => x"23267101",
         281 => x"23248101",
         282 => x"23229101",
         283 => x"2320a101",
         284 => x"130a0500",
         285 => x"93040000",
         286 => x"63dc0500",
         287 => x"b337a000",
         288 => x"b305b040",
         289 => x"b385f540",
         290 => x"330aa040",
         291 => x"9304f0ff",
         292 => x"63dc0600",
         293 => x"b337c000",
         294 => x"b306d040",
         295 => x"93c4f4ff",
         296 => x"b386f640",
         297 => x"3306c040",
         298 => x"930a0600",
         299 => x"93090a00",
         300 => x"13890500",
         301 => x"639a0638",
         302 => x"b7370000",
         303 => x"93874718",
         304 => x"63f6c512",
         305 => x"37070100",
         306 => x"6378e610",
         307 => x"13370610",
         308 => x"13471700",
         309 => x"13173700",
         310 => x"b356e600",
         311 => x"b387d700",
         312 => x"83c70700",
         313 => x"93060002",
         314 => x"b387e700",
         315 => x"3387f640",
         316 => x"638cf600",
         317 => x"3399e500",
         318 => x"b357fa00",
         319 => x"b31ae600",
         320 => x"33e92701",
         321 => x"b319ea00",
         322 => x"13db0a01",
         323 => x"93050b00",
         324 => x"13050900",
         325 => x"939b0a01",
         326 => x"ef108050",
         327 => x"93db0b01",
         328 => x"93050500",
         329 => x"130a0500",
         330 => x"13850b00",
         331 => x"ef10804c",
         332 => x"13040500",
         333 => x"93050b00",
         334 => x"13050900",
         335 => x"ef10c052",
         336 => x"13150501",
         337 => x"13d70901",
         338 => x"3367a700",
         339 => x"13090a00",
         340 => x"637e8700",
         341 => x"33075701",
         342 => x"1309faff",
         343 => x"63685701",
         344 => x"63768700",
         345 => x"1309eaff",
         346 => x"33075701",
         347 => x"33048740",
         348 => x"93050b00",
         349 => x"13050400",
         350 => x"ef10804a",
         351 => x"93050500",
         352 => x"130a0500",
         353 => x"13850b00",
         354 => x"ef10c046",
         355 => x"930b0500",
         356 => x"93050b00",
         357 => x"13050400",
         358 => x"ef10004d",
         359 => x"13970901",
         360 => x"13150501",
         361 => x"13570701",
         362 => x"3367a700",
         363 => x"93060a00",
         364 => x"637c7701",
         365 => x"3387ea00",
         366 => x"9306faff",
         367 => x"63665701",
         368 => x"63747701",
         369 => x"9306eaff",
         370 => x"93170901",
         371 => x"b3e7d700",
         372 => x"13090000",
         373 => x"6f000012",
         374 => x"b7060001",
         375 => x"13070001",
         376 => x"e36cd6ee",
         377 => x"13078001",
         378 => x"6ff01fef",
         379 => x"63140600",
         380 => x"73001000",
         381 => x"37070100",
         382 => x"6378e614",
         383 => x"13370610",
         384 => x"13471700",
         385 => x"13173700",
         386 => x"b356e600",
         387 => x"b387d700",
         388 => x"83c70700",
         389 => x"93060002",
         390 => x"b387e700",
         391 => x"3387f640",
         392 => x"639ef612",
         393 => x"338ac540",
         394 => x"13091000",
         395 => x"93db0a01",
         396 => x"93850b00",
         397 => x"13050a00",
         398 => x"139c0a01",
         399 => x"ef10403e",
         400 => x"135c0c01",
         401 => x"93050500",
         402 => x"930c0500",
         403 => x"13050c00",
         404 => x"ef10403a",
         405 => x"130b0500",
         406 => x"93850b00",
         407 => x"13050a00",
         408 => x"ef108040",
         409 => x"13150501",
         410 => x"13d70901",
         411 => x"3367a700",
         412 => x"138a0c00",
         413 => x"637e6701",
         414 => x"33075701",
         415 => x"138afcff",
         416 => x"63685701",
         417 => x"63766701",
         418 => x"138aecff",
         419 => x"33075701",
         420 => x"33046741",
         421 => x"93850b00",
         422 => x"13050400",
         423 => x"ef104038",
         424 => x"93050500",
         425 => x"130b0500",
         426 => x"13050c00",
         427 => x"ef108034",
         428 => x"130c0500",
         429 => x"93850b00",
         430 => x"13050400",
         431 => x"ef10c03a",
         432 => x"13970901",
         433 => x"13150501",
         434 => x"13570701",
         435 => x"3367a700",
         436 => x"93060b00",
         437 => x"637c8701",
         438 => x"3387ea00",
         439 => x"9306fbff",
         440 => x"63665701",
         441 => x"63748701",
         442 => x"9306ebff",
         443 => x"93170a01",
         444 => x"b3e7d700",
         445 => x"13850700",
         446 => x"93050900",
         447 => x"638a0400",
         448 => x"b337f000",
         449 => x"b3052041",
         450 => x"b385f540",
         451 => x"3305a040",
         452 => x"8320c102",
         453 => x"03248102",
         454 => x"83244102",
         455 => x"03290102",
         456 => x"8329c101",
         457 => x"032a8101",
         458 => x"832a4101",
         459 => x"032b0101",
         460 => x"832bc100",
         461 => x"032c8100",
         462 => x"832c4100",
         463 => x"032d0100",
         464 => x"13010103",
         465 => x"67800000",
         466 => x"b7060001",
         467 => x"13070001",
         468 => x"e36cd6ea",
         469 => x"13078001",
         470 => x"6ff01feb",
         471 => x"b31ae600",
         472 => x"33d9f500",
         473 => x"13dc0a01",
         474 => x"b395e500",
         475 => x"b357fa00",
         476 => x"33ebb700",
         477 => x"b319ea00",
         478 => x"93050c00",
         479 => x"13050900",
         480 => x"139a0a01",
         481 => x"ef10c029",
         482 => x"135a0a01",
         483 => x"93050500",
         484 => x"930b0500",
         485 => x"13050a00",
         486 => x"ef10c025",
         487 => x"13040500",
         488 => x"93050c00",
         489 => x"13050900",
         490 => x"ef10002c",
         491 => x"13150501",
         492 => x"13570b01",
         493 => x"3367a700",
         494 => x"13890b00",
         495 => x"637e8700",
         496 => x"33075701",
         497 => x"1389fbff",
         498 => x"63685701",
         499 => x"63768700",
         500 => x"1389ebff",
         501 => x"33075701",
         502 => x"33048740",
         503 => x"93050c00",
         504 => x"13050400",
         505 => x"ef10c023",
         506 => x"93050500",
         507 => x"930b0500",
         508 => x"13050a00",
         509 => x"ef100020",
         510 => x"130a0500",
         511 => x"93050c00",
         512 => x"13050400",
         513 => x"ef104026",
         514 => x"93170b01",
         515 => x"13150501",
         516 => x"93d70701",
         517 => x"b3e7a700",
         518 => x"13870b00",
         519 => x"63fe4701",
         520 => x"b3875701",
         521 => x"1387fbff",
         522 => x"63e85701",
         523 => x"63f64701",
         524 => x"1387ebff",
         525 => x"b3875701",
         526 => x"13190901",
         527 => x"338a4741",
         528 => x"3369e900",
         529 => x"6ff09fde",
         530 => x"63ecd51e",
         531 => x"b7070100",
         532 => x"63f4f604",
         533 => x"13b50610",
         534 => x"13451500",
         535 => x"13153500",
         536 => x"b7370000",
         537 => x"33d7a600",
         538 => x"93874718",
         539 => x"b387e700",
         540 => x"03c70700",
         541 => x"93070002",
         542 => x"3307a700",
         543 => x"3389e740",
         544 => x"6396e702",
         545 => x"93071000",
         546 => x"e3e6b6e6",
         547 => x"b337ca00",
         548 => x"93c71700",
         549 => x"6ff01fe6",
         550 => x"b7070001",
         551 => x"13050001",
         552 => x"e3e0f6fc",
         553 => x"13058001",
         554 => x"6ff09ffb",
         555 => x"b35be600",
         556 => x"b3962601",
         557 => x"b3ebdb00",
         558 => x"b3dae500",
         559 => x"93dc0b01",
         560 => x"3357ea00",
         561 => x"b3952501",
         562 => x"336bb700",
         563 => x"13850a00",
         564 => x"93850c00",
         565 => x"139c0b01",
         566 => x"33142601",
         567 => x"135c0c01",
         568 => x"ef100014",
         569 => x"93050500",
         570 => x"130d0500",
         571 => x"13050c00",
         572 => x"ef104010",
         573 => x"93090500",
         574 => x"93850c00",
         575 => x"13850a00",
         576 => x"ef108016",
         577 => x"13150501",
         578 => x"13560b01",
         579 => x"3366a600",
         580 => x"930a0d00",
         581 => x"637e3601",
         582 => x"33067601",
         583 => x"930afdff",
         584 => x"63687601",
         585 => x"63763601",
         586 => x"930aedff",
         587 => x"33067601",
         588 => x"b3093641",
         589 => x"93850c00",
         590 => x"13850900",
         591 => x"ef10400e",
         592 => x"93050500",
         593 => x"130d0500",
         594 => x"13050c00",
         595 => x"ef10800a",
         596 => x"130c0500",
         597 => x"93850c00",
         598 => x"13850900",
         599 => x"ef10c010",
         600 => x"13170b01",
         601 => x"13150501",
         602 => x"13570701",
         603 => x"3367a700",
         604 => x"93060d00",
         605 => x"637e8701",
         606 => x"33077701",
         607 => x"9306fdff",
         608 => x"63687701",
         609 => x"63768701",
         610 => x"9306edff",
         611 => x"33077701",
         612 => x"93970a01",
         613 => x"370e0100",
         614 => x"b3e7d700",
         615 => x"1303feff",
         616 => x"33088741",
         617 => x"33f76700",
         618 => x"33736400",
         619 => x"93de0701",
         620 => x"13540401",
         621 => x"13050700",
         622 => x"93050300",
         623 => x"ef108003",
         624 => x"93080500",
         625 => x"93050400",
         626 => x"13050700",
         627 => x"ef108002",
         628 => x"13070500",
         629 => x"93050300",
         630 => x"13850e00",
         631 => x"ef108001",
         632 => x"13030500",
         633 => x"93050400",
         634 => x"13850e00",
         635 => x"ef108000",
         636 => x"33076700",
         637 => x"93d60801",
         638 => x"3307d700",
         639 => x"63746700",
         640 => x"3305c501",
         641 => x"93560701",
         642 => x"b386a600",
         643 => x"6366d802",
         644 => x"e310d8bc",
         645 => x"37060100",
         646 => x"1306f6ff",
         647 => x"3377c700",
         648 => x"13170701",
         649 => x"b3f8c800",
         650 => x"b3162a01",
         651 => x"33071701",
         652 => x"13090000",
         653 => x"e3f0e6cc",
         654 => x"9387f7ff",
         655 => x"6ff05fb9",
         656 => x"13090000",
         657 => x"93070000",
         658 => x"6ff0dfca",
         659 => x"130101fc",
         660 => x"232a9102",
         661 => x"232e1102",
         662 => x"232c8102",
         663 => x"23282103",
         664 => x"23263103",
         665 => x"23244103",
         666 => x"23225103",
         667 => x"23206103",
         668 => x"232e7101",
         669 => x"232c8101",
         670 => x"232a9101",
         671 => x"2328a101",
         672 => x"2326b101",
         673 => x"93040000",
         674 => x"63dc0500",
         675 => x"b337a000",
         676 => x"b305b040",
         677 => x"b385f540",
         678 => x"3305a040",
         679 => x"9304f0ff",
         680 => x"63da0600",
         681 => x"b337c000",
         682 => x"b306d040",
         683 => x"b386f640",
         684 => x"3306c040",
         685 => x"130a0600",
         686 => x"13040500",
         687 => x"13890500",
         688 => x"63960626",
         689 => x"b7370000",
         690 => x"93874718",
         691 => x"63fac514",
         692 => x"37070100",
         693 => x"637ce612",
         694 => x"13370610",
         695 => x"13471700",
         696 => x"13173700",
         697 => x"b356e600",
         698 => x"b387d700",
         699 => x"83c70700",
         700 => x"b387e700",
         701 => x"13070002",
         702 => x"b309f740",
         703 => x"630cf700",
         704 => x"b3953501",
         705 => x"b357f500",
         706 => x"331a3601",
         707 => x"33e9b700",
         708 => x"33143501",
         709 => x"135b0a01",
         710 => x"93050b00",
         711 => x"931b0a01",
         712 => x"13050900",
         713 => x"ef00d06f",
         714 => x"93db0b01",
         715 => x"93850b00",
         716 => x"ef00506c",
         717 => x"930a0500",
         718 => x"93050b00",
         719 => x"13050900",
         720 => x"ef009072",
         721 => x"13150501",
         722 => x"93570401",
         723 => x"b3e7a700",
         724 => x"63fa5701",
         725 => x"b3874701",
         726 => x"63e64701",
         727 => x"63f45701",
         728 => x"b3874701",
         729 => x"33895741",
         730 => x"93050b00",
         731 => x"13050900",
         732 => x"ef00106b",
         733 => x"93850b00",
         734 => x"ef00d067",
         735 => x"930a0500",
         736 => x"93050b00",
         737 => x"13050900",
         738 => x"ef00106e",
         739 => x"13140401",
         740 => x"13150501",
         741 => x"13540401",
         742 => x"3364a400",
         743 => x"637a5401",
         744 => x"33044401",
         745 => x"63664401",
         746 => x"63745401",
         747 => x"33044401",
         748 => x"33045441",
         749 => x"33553401",
         750 => x"93050000",
         751 => x"638a0400",
         752 => x"b337a000",
         753 => x"b305b040",
         754 => x"b385f540",
         755 => x"3305a040",
         756 => x"8320c103",
         757 => x"03248103",
         758 => x"83244103",
         759 => x"03290103",
         760 => x"8329c102",
         761 => x"032a8102",
         762 => x"832a4102",
         763 => x"032b0102",
         764 => x"832bc101",
         765 => x"032c8101",
         766 => x"832c4101",
         767 => x"032d0101",
         768 => x"832dc100",
         769 => x"13010104",
         770 => x"67800000",
         771 => x"b7060001",
         772 => x"13070001",
         773 => x"e368d6ec",
         774 => x"13078001",
         775 => x"6ff09fec",
         776 => x"63140600",
         777 => x"73001000",
         778 => x"37070100",
         779 => x"6376e60e",
         780 => x"13370610",
         781 => x"13471700",
         782 => x"13173700",
         783 => x"b356e600",
         784 => x"b387d700",
         785 => x"83c70700",
         786 => x"3389c540",
         787 => x"b387e700",
         788 => x"13070002",
         789 => x"b309f740",
         790 => x"e30ef7ea",
         791 => x"331a3601",
         792 => x"33dcf500",
         793 => x"935b0a01",
         794 => x"b357f500",
         795 => x"b3953501",
         796 => x"b3eab700",
         797 => x"33143501",
         798 => x"93850b00",
         799 => x"131b0a01",
         800 => x"13050c00",
         801 => x"ef00d059",
         802 => x"135b0b01",
         803 => x"93050b00",
         804 => x"ef005056",
         805 => x"13090500",
         806 => x"93850b00",
         807 => x"13050c00",
         808 => x"ef00905c",
         809 => x"13150501",
         810 => x"13d70a01",
         811 => x"3367a700",
         812 => x"637a2701",
         813 => x"33074701",
         814 => x"63664701",
         815 => x"63742701",
         816 => x"33074701",
         817 => x"33092741",
         818 => x"93850b00",
         819 => x"13050900",
         820 => x"ef001055",
         821 => x"93050b00",
         822 => x"ef00d051",
         823 => x"130b0500",
         824 => x"93850b00",
         825 => x"13050900",
         826 => x"ef001058",
         827 => x"93970a01",
         828 => x"13150501",
         829 => x"93d70701",
         830 => x"b3e7a700",
         831 => x"63fa6701",
         832 => x"b3874701",
         833 => x"63e64701",
         834 => x"63f46701",
         835 => x"b3874701",
         836 => x"33896741",
         837 => x"6ff01fe0",
         838 => x"b7060001",
         839 => x"13070001",
         840 => x"e36ed6f0",
         841 => x"13078001",
         842 => x"6ff05ff1",
         843 => x"e3e8d5e8",
         844 => x"b7070100",
         845 => x"63fef604",
         846 => x"93b70610",
         847 => x"93c71700",
         848 => x"93973700",
         849 => x"37370000",
         850 => x"33d8f600",
         851 => x"13074718",
         852 => x"33070701",
         853 => x"034a0700",
         854 => x"330afa00",
         855 => x"93070002",
         856 => x"b3894741",
         857 => x"63904705",
         858 => x"63e4b600",
         859 => x"636cc500",
         860 => x"3306c540",
         861 => x"b386d540",
         862 => x"b335c500",
         863 => x"3389b640",
         864 => x"13040600",
         865 => x"13050400",
         866 => x"93050900",
         867 => x"6ff01fe3",
         868 => x"37070001",
         869 => x"93070001",
         870 => x"e3e6e6fa",
         871 => x"93078001",
         872 => x"6ff05ffa",
         873 => x"b3963601",
         874 => x"b35b4601",
         875 => x"b3ebdb00",
         876 => x"33dd4501",
         877 => x"33544501",
         878 => x"b3953501",
         879 => x"13dc0b01",
         880 => x"3364b400",
         881 => x"33193501",
         882 => x"93050c00",
         883 => x"13050d00",
         884 => x"939c0b01",
         885 => x"b31a3601",
         886 => x"93dc0c01",
         887 => x"ef005044",
         888 => x"93050500",
         889 => x"930d0500",
         890 => x"13850c00",
         891 => x"ef009040",
         892 => x"130b0500",
         893 => x"93050c00",
         894 => x"13050d00",
         895 => x"ef00d046",
         896 => x"13150501",
         897 => x"93570401",
         898 => x"b3e7a700",
         899 => x"138d0d00",
         900 => x"63fe6701",
         901 => x"b3877701",
         902 => x"138dfdff",
         903 => x"63e87701",
         904 => x"63f66701",
         905 => x"138dedff",
         906 => x"b3877701",
         907 => x"338b6741",
         908 => x"93050c00",
         909 => x"13050b00",
         910 => x"ef00903e",
         911 => x"93050500",
         912 => x"930d0500",
         913 => x"13850c00",
         914 => x"ef00d03a",
         915 => x"93050c00",
         916 => x"930c0500",
         917 => x"13050b00",
         918 => x"ef001041",
         919 => x"93150401",
         920 => x"13150501",
         921 => x"93d50501",
         922 => x"b3e5a500",
         923 => x"13870d00",
         924 => x"63fe9501",
         925 => x"b3857501",
         926 => x"1387fdff",
         927 => x"63e87501",
         928 => x"63f69501",
         929 => x"1387edff",
         930 => x"b3857501",
         931 => x"37030100",
         932 => x"131d0d01",
         933 => x"336ded00",
         934 => x"1307f3ff",
         935 => x"337eed00",
         936 => x"33f7ea00",
         937 => x"b3879541",
         938 => x"135d0d01",
         939 => x"93d80a01",
         940 => x"13050e00",
         941 => x"93050700",
         942 => x"ef00d033",
         943 => x"13080500",
         944 => x"93850800",
         945 => x"13050e00",
         946 => x"ef00d032",
         947 => x"13040500",
         948 => x"93050700",
         949 => x"13050d00",
         950 => x"ef00d031",
         951 => x"13070500",
         952 => x"93850800",
         953 => x"13050d00",
         954 => x"ef00d030",
         955 => x"3304e400",
         956 => x"93560801",
         957 => x"3304d400",
         958 => x"6374e400",
         959 => x"33056500",
         960 => x"b7060100",
         961 => x"9386f6ff",
         962 => x"13570401",
         963 => x"3374d400",
         964 => x"13140401",
         965 => x"3378d800",
         966 => x"3307a700",
         967 => x"33040401",
         968 => x"63e6e700",
         969 => x"639ee700",
         970 => x"637c8900",
         971 => x"33065441",
         972 => x"3334c400",
         973 => x"33047401",
         974 => x"33078740",
         975 => x"13040600",
         976 => x"33048940",
         977 => x"33398900",
         978 => x"b385e740",
         979 => x"b3852541",
         980 => x"339a4501",
         981 => x"33543401",
         982 => x"33658a00",
         983 => x"b3d53501",
         984 => x"6ff0dfc5",
         985 => x"130101fd",
         986 => x"232e3101",
         987 => x"23261102",
         988 => x"23248102",
         989 => x"23229102",
         990 => x"23202103",
         991 => x"232c4101",
         992 => x"232a5101",
         993 => x"23286101",
         994 => x"23267101",
         995 => x"23248101",
         996 => x"23229101",
         997 => x"93090500",
         998 => x"63940638",
         999 => x"b7370000",
        1000 => x"130a0600",
        1001 => x"93040500",
        1002 => x"93874718",
        1003 => x"63f8c512",
        1004 => x"37070100",
        1005 => x"13890500",
        1006 => x"6378e610",
        1007 => x"13370610",
        1008 => x"13471700",
        1009 => x"13173700",
        1010 => x"b356e600",
        1011 => x"b387d700",
        1012 => x"83c70700",
        1013 => x"93060002",
        1014 => x"b387e700",
        1015 => x"3387f640",
        1016 => x"638cf600",
        1017 => x"3399e500",
        1018 => x"b3d7f900",
        1019 => x"331ae600",
        1020 => x"33e92701",
        1021 => x"b394e900",
        1022 => x"935a0a01",
        1023 => x"93850a00",
        1024 => x"13050900",
        1025 => x"131b0a01",
        1026 => x"ef009021",
        1027 => x"135b0b01",
        1028 => x"93050500",
        1029 => x"93090500",
        1030 => x"13050b00",
        1031 => x"ef00901d",
        1032 => x"13040500",
        1033 => x"93850a00",
        1034 => x"13050900",
        1035 => x"ef00d023",
        1036 => x"13150501",
        1037 => x"13d70401",
        1038 => x"3367a700",
        1039 => x"13890900",
        1040 => x"637e8700",
        1041 => x"33074701",
        1042 => x"1389f9ff",
        1043 => x"63684701",
        1044 => x"63768700",
        1045 => x"1389e9ff",
        1046 => x"33074701",
        1047 => x"33048740",
        1048 => x"93850a00",
        1049 => x"13050400",
        1050 => x"ef00901b",
        1051 => x"93050500",
        1052 => x"93090500",
        1053 => x"13050b00",
        1054 => x"ef00d017",
        1055 => x"130b0500",
        1056 => x"93850a00",
        1057 => x"13050400",
        1058 => x"ef00101e",
        1059 => x"13970401",
        1060 => x"13150501",
        1061 => x"13570701",
        1062 => x"3367a700",
        1063 => x"93860900",
        1064 => x"637c6701",
        1065 => x"3307ea00",
        1066 => x"9386f9ff",
        1067 => x"63664701",
        1068 => x"63746701",
        1069 => x"9386e9ff",
        1070 => x"93170901",
        1071 => x"b3e7d700",
        1072 => x"13090000",
        1073 => x"6f000012",
        1074 => x"b7060001",
        1075 => x"13070001",
        1076 => x"e36cd6ee",
        1077 => x"13078001",
        1078 => x"6ff01fef",
        1079 => x"63140600",
        1080 => x"73001000",
        1081 => x"37070100",
        1082 => x"637ce612",
        1083 => x"13370610",
        1084 => x"13471700",
        1085 => x"13173700",
        1086 => x"b356e600",
        1087 => x"b387d700",
        1088 => x"83c70700",
        1089 => x"93060002",
        1090 => x"b387e700",
        1091 => x"3387f640",
        1092 => x"6392f612",
        1093 => x"b389c540",
        1094 => x"13091000",
        1095 => x"135b0a01",
        1096 => x"93050b00",
        1097 => x"13850900",
        1098 => x"931b0a01",
        1099 => x"ef00500f",
        1100 => x"93db0b01",
        1101 => x"93050500",
        1102 => x"130c0500",
        1103 => x"13850b00",
        1104 => x"ef00500b",
        1105 => x"930a0500",
        1106 => x"93050b00",
        1107 => x"13850900",
        1108 => x"ef009011",
        1109 => x"13150501",
        1110 => x"13d70401",
        1111 => x"3367a700",
        1112 => x"93090c00",
        1113 => x"637e5701",
        1114 => x"33074701",
        1115 => x"9309fcff",
        1116 => x"63684701",
        1117 => x"63765701",
        1118 => x"9309ecff",
        1119 => x"33074701",
        1120 => x"33045741",
        1121 => x"93050b00",
        1122 => x"13050400",
        1123 => x"ef005009",
        1124 => x"93050500",
        1125 => x"930a0500",
        1126 => x"13850b00",
        1127 => x"ef009005",
        1128 => x"930b0500",
        1129 => x"93050b00",
        1130 => x"13050400",
        1131 => x"ef00d00b",
        1132 => x"13970401",
        1133 => x"13150501",
        1134 => x"13570701",
        1135 => x"3367a700",
        1136 => x"93860a00",
        1137 => x"637c7701",
        1138 => x"3307ea00",
        1139 => x"9386faff",
        1140 => x"63664701",
        1141 => x"63747701",
        1142 => x"9386eaff",
        1143 => x"93970901",
        1144 => x"b3e7d700",
        1145 => x"8320c102",
        1146 => x"03248102",
        1147 => x"83244102",
        1148 => x"8329c101",
        1149 => x"032a8101",
        1150 => x"832a4101",
        1151 => x"032b0101",
        1152 => x"832bc100",
        1153 => x"032c8100",
        1154 => x"832c4100",
        1155 => x"93050900",
        1156 => x"13850700",
        1157 => x"03290102",
        1158 => x"13010103",
        1159 => x"67800000",
        1160 => x"b7060001",
        1161 => x"13070001",
        1162 => x"e368d6ec",
        1163 => x"13078001",
        1164 => x"6ff09fec",
        1165 => x"331ae600",
        1166 => x"33d9f500",
        1167 => x"935b0a01",
        1168 => x"b395e500",
        1169 => x"b3d7f900",
        1170 => x"b3eab700",
        1171 => x"b394e900",
        1172 => x"93850b00",
        1173 => x"13050900",
        1174 => x"93190a01",
        1175 => x"ef00407c",
        1176 => x"93d90901",
        1177 => x"93050500",
        1178 => x"130b0500",
        1179 => x"13850900",
        1180 => x"ef004078",
        1181 => x"13040500",
        1182 => x"93850b00",
        1183 => x"13050900",
        1184 => x"ef00807e",
        1185 => x"13150501",
        1186 => x"13d70a01",
        1187 => x"3367a700",
        1188 => x"13090b00",
        1189 => x"637e8700",
        1190 => x"33074701",
        1191 => x"1309fbff",
        1192 => x"63684701",
        1193 => x"63768700",
        1194 => x"1309ebff",
        1195 => x"33074701",
        1196 => x"33048740",
        1197 => x"93850b00",
        1198 => x"13050400",
        1199 => x"ef004076",
        1200 => x"93050500",
        1201 => x"130b0500",
        1202 => x"13850900",
        1203 => x"ef008072",
        1204 => x"93090500",
        1205 => x"93850b00",
        1206 => x"13050400",
        1207 => x"ef00c078",
        1208 => x"93970a01",
        1209 => x"13150501",
        1210 => x"93d70701",
        1211 => x"b3e7a700",
        1212 => x"13070b00",
        1213 => x"63fe3701",
        1214 => x"b3874701",
        1215 => x"1307fbff",
        1216 => x"63e84701",
        1217 => x"63f63701",
        1218 => x"1307ebff",
        1219 => x"b3874701",
        1220 => x"13190901",
        1221 => x"b3893741",
        1222 => x"3369e900",
        1223 => x"6ff01fe0",
        1224 => x"63ecd51e",
        1225 => x"b7070100",
        1226 => x"63f4f604",
        1227 => x"13b50610",
        1228 => x"13451500",
        1229 => x"13153500",
        1230 => x"b7370000",
        1231 => x"33d7a600",
        1232 => x"93874718",
        1233 => x"b387e700",
        1234 => x"03c70700",
        1235 => x"93070002",
        1236 => x"3307a700",
        1237 => x"3389e740",
        1238 => x"6396e702",
        1239 => x"93071000",
        1240 => x"e3e2b6e8",
        1241 => x"b3b7c900",
        1242 => x"93c71700",
        1243 => x"6ff09fe7",
        1244 => x"b7070001",
        1245 => x"13050001",
        1246 => x"e3e0f6fc",
        1247 => x"13058001",
        1248 => x"6ff09ffb",
        1249 => x"b3962601",
        1250 => x"335be600",
        1251 => x"336bdb00",
        1252 => x"33dae500",
        1253 => x"135c0b01",
        1254 => x"33d7e900",
        1255 => x"b3952501",
        1256 => x"b36ab700",
        1257 => x"13050a00",
        1258 => x"93050c00",
        1259 => x"931b0b01",
        1260 => x"b3142601",
        1261 => x"93db0b01",
        1262 => x"ef008066",
        1263 => x"93050500",
        1264 => x"930c0500",
        1265 => x"13850b00",
        1266 => x"ef00c062",
        1267 => x"13040500",
        1268 => x"93050c00",
        1269 => x"13050a00",
        1270 => x"ef000069",
        1271 => x"13150501",
        1272 => x"93d60a01",
        1273 => x"b3e6a600",
        1274 => x"138a0c00",
        1275 => x"63fe8600",
        1276 => x"b3866601",
        1277 => x"138afcff",
        1278 => x"63e86601",
        1279 => x"63f68600",
        1280 => x"138aecff",
        1281 => x"b3866601",
        1282 => x"33848640",
        1283 => x"93050c00",
        1284 => x"13050400",
        1285 => x"ef00c060",
        1286 => x"93050500",
        1287 => x"930c0500",
        1288 => x"13850b00",
        1289 => x"ef00005d",
        1290 => x"930b0500",
        1291 => x"93050c00",
        1292 => x"13050400",
        1293 => x"ef004063",
        1294 => x"13970a01",
        1295 => x"13150501",
        1296 => x"13570701",
        1297 => x"3367a700",
        1298 => x"93860c00",
        1299 => x"637e7701",
        1300 => x"33076701",
        1301 => x"9386fcff",
        1302 => x"63686701",
        1303 => x"63767701",
        1304 => x"9386ecff",
        1305 => x"33076701",
        1306 => x"93170a01",
        1307 => x"370e0100",
        1308 => x"b3e7d700",
        1309 => x"1303feff",
        1310 => x"33087741",
        1311 => x"33f76700",
        1312 => x"33f36400",
        1313 => x"93de0701",
        1314 => x"93d40401",
        1315 => x"13050700",
        1316 => x"93050300",
        1317 => x"ef000056",
        1318 => x"93080500",
        1319 => x"93850400",
        1320 => x"13050700",
        1321 => x"ef000055",
        1322 => x"13070500",
        1323 => x"93050300",
        1324 => x"13850e00",
        1325 => x"ef000054",
        1326 => x"13030500",
        1327 => x"93850400",
        1328 => x"13850e00",
        1329 => x"ef000053",
        1330 => x"33076700",
        1331 => x"93d60801",
        1332 => x"3307d700",
        1333 => x"63746700",
        1334 => x"3305c501",
        1335 => x"93560701",
        1336 => x"b386a600",
        1337 => x"6366d802",
        1338 => x"e31cd8bc",
        1339 => x"37060100",
        1340 => x"1306f6ff",
        1341 => x"3377c700",
        1342 => x"13170701",
        1343 => x"b3f8c800",
        1344 => x"b3962901",
        1345 => x"33071701",
        1346 => x"13090000",
        1347 => x"e3fce6cc",
        1348 => x"9387f7ff",
        1349 => x"6ff0dfba",
        1350 => x"13090000",
        1351 => x"93070000",
        1352 => x"6ff05fcc",
        1353 => x"130101fd",
        1354 => x"23248102",
        1355 => x"23229102",
        1356 => x"23261102",
        1357 => x"23202103",
        1358 => x"232e3101",
        1359 => x"232c4101",
        1360 => x"232a5101",
        1361 => x"23286101",
        1362 => x"23267101",
        1363 => x"23248101",
        1364 => x"23229101",
        1365 => x"2320a101",
        1366 => x"13040500",
        1367 => x"93840500",
        1368 => x"639c0624",
        1369 => x"b7370000",
        1370 => x"130a0600",
        1371 => x"93874718",
        1372 => x"63fec512",
        1373 => x"37070100",
        1374 => x"6370e612",
        1375 => x"13370610",
        1376 => x"13471700",
        1377 => x"13173700",
        1378 => x"b356e600",
        1379 => x"b387d700",
        1380 => x"83c70700",
        1381 => x"b387e700",
        1382 => x"13070002",
        1383 => x"3309f740",
        1384 => x"630cf700",
        1385 => x"b3952501",
        1386 => x"b357f500",
        1387 => x"331a2601",
        1388 => x"b3e4b700",
        1389 => x"33142501",
        1390 => x"935a0a01",
        1391 => x"93850a00",
        1392 => x"131b0a01",
        1393 => x"13850400",
        1394 => x"ef008045",
        1395 => x"135b0b01",
        1396 => x"93050b00",
        1397 => x"ef000042",
        1398 => x"93090500",
        1399 => x"93850a00",
        1400 => x"13850400",
        1401 => x"ef004048",
        1402 => x"13150501",
        1403 => x"93570401",
        1404 => x"b3e7a700",
        1405 => x"63fa3701",
        1406 => x"b3874701",
        1407 => x"63e64701",
        1408 => x"63f43701",
        1409 => x"b3874701",
        1410 => x"b3843741",
        1411 => x"93850a00",
        1412 => x"13850400",
        1413 => x"ef00c040",
        1414 => x"93050b00",
        1415 => x"ef00803d",
        1416 => x"93090500",
        1417 => x"93850a00",
        1418 => x"13850400",
        1419 => x"ef00c043",
        1420 => x"13140401",
        1421 => x"13150501",
        1422 => x"13540401",
        1423 => x"3364a400",
        1424 => x"637a3401",
        1425 => x"33044401",
        1426 => x"63664401",
        1427 => x"63743401",
        1428 => x"33044401",
        1429 => x"33043441",
        1430 => x"33552401",
        1431 => x"93050000",
        1432 => x"8320c102",
        1433 => x"03248102",
        1434 => x"83244102",
        1435 => x"03290102",
        1436 => x"8329c101",
        1437 => x"032a8101",
        1438 => x"832a4101",
        1439 => x"032b0101",
        1440 => x"832bc100",
        1441 => x"032c8100",
        1442 => x"832c4100",
        1443 => x"032d0100",
        1444 => x"13010103",
        1445 => x"67800000",
        1446 => x"b7060001",
        1447 => x"13070001",
        1448 => x"e364d6ee",
        1449 => x"13078001",
        1450 => x"6ff01fee",
        1451 => x"63140600",
        1452 => x"73001000",
        1453 => x"37070100",
        1454 => x"6376e60e",
        1455 => x"13370610",
        1456 => x"13471700",
        1457 => x"13173700",
        1458 => x"b356e600",
        1459 => x"b387d700",
        1460 => x"83c70700",
        1461 => x"b384c540",
        1462 => x"b387e700",
        1463 => x"13070002",
        1464 => x"3309f740",
        1465 => x"e30af7ec",
        1466 => x"331a2601",
        1467 => x"b3dbf500",
        1468 => x"135b0a01",
        1469 => x"b357f500",
        1470 => x"b3952501",
        1471 => x"b3e9b700",
        1472 => x"33142501",
        1473 => x"93050b00",
        1474 => x"931a0a01",
        1475 => x"13850b00",
        1476 => x"ef000031",
        1477 => x"93da0a01",
        1478 => x"93850a00",
        1479 => x"ef00802d",
        1480 => x"93040500",
        1481 => x"93050b00",
        1482 => x"13850b00",
        1483 => x"ef00c033",
        1484 => x"13150501",
        1485 => x"13d70901",
        1486 => x"3367a700",
        1487 => x"637a9700",
        1488 => x"33074701",
        1489 => x"63664701",
        1490 => x"63749700",
        1491 => x"33074701",
        1492 => x"b3049740",
        1493 => x"93050b00",
        1494 => x"13850400",
        1495 => x"ef00402c",
        1496 => x"93850a00",
        1497 => x"ef000029",
        1498 => x"930a0500",
        1499 => x"93050b00",
        1500 => x"13850400",
        1501 => x"ef00402f",
        1502 => x"93970901",
        1503 => x"13150501",
        1504 => x"93d70701",
        1505 => x"b3e7a700",
        1506 => x"63fa5701",
        1507 => x"b3874701",
        1508 => x"63e64701",
        1509 => x"63f45701",
        1510 => x"b3874701",
        1511 => x"b3845741",
        1512 => x"6ff09fe1",
        1513 => x"b7060001",
        1514 => x"13070001",
        1515 => x"e36ed6f0",
        1516 => x"13078001",
        1517 => x"6ff05ff1",
        1518 => x"e3e4d5ea",
        1519 => x"b7070100",
        1520 => x"63fef604",
        1521 => x"93b70610",
        1522 => x"93c71700",
        1523 => x"93973700",
        1524 => x"37370000",
        1525 => x"33d8f600",
        1526 => x"13074718",
        1527 => x"33070701",
        1528 => x"83490700",
        1529 => x"b389f900",
        1530 => x"93070002",
        1531 => x"33893741",
        1532 => x"63903705",
        1533 => x"63e4b600",
        1534 => x"636cc500",
        1535 => x"3306c540",
        1536 => x"b386d540",
        1537 => x"b335c500",
        1538 => x"b384b640",
        1539 => x"13040600",
        1540 => x"13050400",
        1541 => x"93850400",
        1542 => x"6ff09fe4",
        1543 => x"37070001",
        1544 => x"93070001",
        1545 => x"e3e6e6fa",
        1546 => x"93078001",
        1547 => x"6ff05ffa",
        1548 => x"b3962601",
        1549 => x"335b3601",
        1550 => x"336bdb00",
        1551 => x"b3d43501",
        1552 => x"335a3501",
        1553 => x"b3952501",
        1554 => x"935c0b01",
        1555 => x"336aba00",
        1556 => x"b31a2501",
        1557 => x"93850c00",
        1558 => x"13850400",
        1559 => x"131c0b01",
        1560 => x"b31b2601",
        1561 => x"135c0c01",
        1562 => x"ef00801b",
        1563 => x"93050500",
        1564 => x"130d0500",
        1565 => x"13050c00",
        1566 => x"ef00c017",
        1567 => x"13040500",
        1568 => x"93850c00",
        1569 => x"13850400",
        1570 => x"ef00001e",
        1571 => x"13150501",
        1572 => x"93570a01",
        1573 => x"b3e7a700",
        1574 => x"93040d00",
        1575 => x"63fe8700",
        1576 => x"b3876701",
        1577 => x"9304fdff",
        1578 => x"63e86701",
        1579 => x"63f68700",
        1580 => x"9304edff",
        1581 => x"b3876701",
        1582 => x"33848740",
        1583 => x"93850c00",
        1584 => x"13050400",
        1585 => x"ef00c015",
        1586 => x"93050500",
        1587 => x"130d0500",
        1588 => x"13050c00",
        1589 => x"ef000012",
        1590 => x"93850c00",
        1591 => x"130c0500",
        1592 => x"13050400",
        1593 => x"ef004018",
        1594 => x"93150a01",
        1595 => x"13150501",
        1596 => x"93d50501",
        1597 => x"b3e5a500",
        1598 => x"93070d00",
        1599 => x"63fe8501",
        1600 => x"b3856501",
        1601 => x"9307fdff",
        1602 => x"63e86501",
        1603 => x"63f68501",
        1604 => x"9307edff",
        1605 => x"b3856501",
        1606 => x"b70e0100",
        1607 => x"93940401",
        1608 => x"b3e4f400",
        1609 => x"9387feff",
        1610 => x"b3f8f400",
        1611 => x"b3f7fb00",
        1612 => x"33878541",
        1613 => x"93d40401",
        1614 => x"13de0b01",
        1615 => x"13850800",
        1616 => x"93850700",
        1617 => x"ef00000b",
        1618 => x"13080500",
        1619 => x"93050e00",
        1620 => x"13850800",
        1621 => x"ef00000a",
        1622 => x"93080500",
        1623 => x"93850700",
        1624 => x"13850400",
        1625 => x"ef000009",
        1626 => x"13030500",
        1627 => x"93050e00",
        1628 => x"13850400",
        1629 => x"ef000008",
        1630 => x"93570801",
        1631 => x"b3886800",
        1632 => x"b3871701",
        1633 => x"13060500",
        1634 => x"63f46700",
        1635 => x"3306d501",
        1636 => x"93d60701",
        1637 => x"b386c600",
        1638 => x"37060100",
        1639 => x"1306f6ff",
        1640 => x"b3f7c700",
        1641 => x"93970701",
        1642 => x"3378c800",
        1643 => x"b3870701",
        1644 => x"6366d700",
        1645 => x"631ed700",
        1646 => x"63fcfa00",
        1647 => x"33867741",
        1648 => x"b3b7c700",
        1649 => x"b3876701",
        1650 => x"b386f640",
        1651 => x"93070600",
        1652 => x"b387fa40",
        1653 => x"b3bafa00",
        1654 => x"b305d740",
        1655 => x"b3855541",
        1656 => x"b3993501",
        1657 => x"b3d72701",
        1658 => x"33e5f900",
        1659 => x"b3d52501",
        1660 => x"6ff01fc7",
        1661 => x"13060500",
        1662 => x"13050000",
        1663 => x"93f61500",
        1664 => x"63840600",
        1665 => x"3305c500",
        1666 => x"93d51500",
        1667 => x"13161600",
        1668 => x"e39605fe",
        1669 => x"67800000",
        1670 => x"63400506",
        1671 => x"63c60506",
        1672 => x"13860500",
        1673 => x"93050500",
        1674 => x"1305f0ff",
        1675 => x"630c0602",
        1676 => x"93061000",
        1677 => x"637ab600",
        1678 => x"6358c000",
        1679 => x"13161600",
        1680 => x"93961600",
        1681 => x"e36ab6fe",
        1682 => x"13050000",
        1683 => x"63e6c500",
        1684 => x"b385c540",
        1685 => x"3365d500",
        1686 => x"93d61600",
        1687 => x"13561600",
        1688 => x"e39606fe",
        1689 => x"67800000",
        1690 => x"93820000",
        1691 => x"eff05ffb",
        1692 => x"13850500",
        1693 => x"67800200",
        1694 => x"3305a040",
        1695 => x"6348b000",
        1696 => x"b305b040",
        1697 => x"6ff0dff9",
        1698 => x"b305b040",
        1699 => x"93820000",
        1700 => x"eff01ff9",
        1701 => x"3305a040",
        1702 => x"67800200",
        1703 => x"93820000",
        1704 => x"63ca0500",
        1705 => x"634c0500",
        1706 => x"eff09ff7",
        1707 => x"13850500",
        1708 => x"67800200",
        1709 => x"b305b040",
        1710 => x"e35805fe",
        1711 => x"3305a040",
        1712 => x"eff01ff6",
        1713 => x"3305b040",
        1714 => x"67800200",
        1715 => x"13030500",
        1716 => x"630a0600",
        1717 => x"2300b300",
        1718 => x"1306f6ff",
        1719 => x"13031300",
        1720 => x"e31a06fe",
        1721 => x"67800000",
        1722 => x"13030500",
        1723 => x"630e0600",
        1724 => x"83830500",
        1725 => x"23007300",
        1726 => x"1306f6ff",
        1727 => x"13031300",
        1728 => x"93851500",
        1729 => x"e31606fe",
        1730 => x"67800000",
        1731 => x"630c0602",
        1732 => x"13030500",
        1733 => x"93061000",
        1734 => x"636ab500",
        1735 => x"9306f0ff",
        1736 => x"1307f6ff",
        1737 => x"3303e300",
        1738 => x"b385e500",
        1739 => x"83830500",
        1740 => x"23007300",
        1741 => x"1306f6ff",
        1742 => x"3303d300",
        1743 => x"b385d500",
        1744 => x"e31606fe",
        1745 => x"67800000",
        1746 => x"03a50186",
        1747 => x"67800000",
        1748 => x"130101ff",
        1749 => x"23248100",
        1750 => x"23261100",
        1751 => x"93070000",
        1752 => x"13040500",
        1753 => x"63880700",
        1754 => x"93050000",
        1755 => x"97000000",
        1756 => x"e7000000",
        1757 => x"b7370000",
        1758 => x"03a58731",
        1759 => x"83278502",
        1760 => x"63840700",
        1761 => x"e7800700",
        1762 => x"13050400",
        1763 => x"ef10c03e",
        1764 => x"130101ff",
        1765 => x"23248100",
        1766 => x"23229100",
        1767 => x"37340000",
        1768 => x"b7340000",
        1769 => x"9387c431",
        1770 => x"1304c431",
        1771 => x"3304f440",
        1772 => x"23202101",
        1773 => x"23261100",
        1774 => x"13542440",
        1775 => x"9384c431",
        1776 => x"13090000",
        1777 => x"63108904",
        1778 => x"b7340000",
        1779 => x"37340000",
        1780 => x"9387c431",
        1781 => x"1304c431",
        1782 => x"3304f440",
        1783 => x"13542440",
        1784 => x"9384c431",
        1785 => x"13090000",
        1786 => x"63188902",
        1787 => x"8320c100",
        1788 => x"03248100",
        1789 => x"83244100",
        1790 => x"03290100",
        1791 => x"13010101",
        1792 => x"67800000",
        1793 => x"83a70400",
        1794 => x"13091900",
        1795 => x"93844400",
        1796 => x"e7800700",
        1797 => x"6ff01ffb",
        1798 => x"83a70400",
        1799 => x"13091900",
        1800 => x"93844400",
        1801 => x"e7800700",
        1802 => x"6ff01ffc",
        1803 => x"130101f7",
        1804 => x"232c8106",
        1805 => x"232a9106",
        1806 => x"232e1106",
        1807 => x"23282107",
        1808 => x"2320e108",
        1809 => x"2322f108",
        1810 => x"23240109",
        1811 => x"23261109",
        1812 => x"93040500",
        1813 => x"13040600",
        1814 => x"63540602",
        1815 => x"9307b008",
        1816 => x"2320f500",
        1817 => x"1305f0ff",
        1818 => x"8320c107",
        1819 => x"03248107",
        1820 => x"83244107",
        1821 => x"03290107",
        1822 => x"13010109",
        1823 => x"67800000",
        1824 => x"93078020",
        1825 => x"231af100",
        1826 => x"2324b100",
        1827 => x"232cb100",
        1828 => x"13860600",
        1829 => x"93070000",
        1830 => x"63040400",
        1831 => x"9307f4ff",
        1832 => x"1309f0ff",
        1833 => x"93060108",
        1834 => x"93058100",
        1835 => x"13850400",
        1836 => x"2328f100",
        1837 => x"232ef100",
        1838 => x"231b2101",
        1839 => x"2322d100",
        1840 => x"ef004045",
        1841 => x"63562501",
        1842 => x"9307b008",
        1843 => x"23a0f400",
        1844 => x"e30c04f8",
        1845 => x"83278100",
        1846 => x"23800700",
        1847 => x"6ff0dff8",
        1848 => x"130101f6",
        1849 => x"232a9106",
        1850 => x"232af108",
        1851 => x"232e1106",
        1852 => x"232c8106",
        1853 => x"23282107",
        1854 => x"2326d108",
        1855 => x"2328e108",
        1856 => x"232c0109",
        1857 => x"232e1109",
        1858 => x"83a40186",
        1859 => x"63d40502",
        1860 => x"9307b008",
        1861 => x"23a0f400",
        1862 => x"1305f0ff",
        1863 => x"8320c107",
        1864 => x"03248107",
        1865 => x"83244107",
        1866 => x"03290107",
        1867 => x"1301010a",
        1868 => x"67800000",
        1869 => x"93078020",
        1870 => x"231af100",
        1871 => x"2324a100",
        1872 => x"232ca100",
        1873 => x"13840500",
        1874 => x"93070000",
        1875 => x"63840500",
        1876 => x"9387f5ff",
        1877 => x"1309f0ff",
        1878 => x"9306c108",
        1879 => x"93058100",
        1880 => x"13850400",
        1881 => x"2328f100",
        1882 => x"232ef100",
        1883 => x"231b2101",
        1884 => x"2322d100",
        1885 => x"ef00003a",
        1886 => x"63562501",
        1887 => x"9307b008",
        1888 => x"23a0f400",
        1889 => x"e30c04f8",
        1890 => x"83278100",
        1891 => x"23800700",
        1892 => x"6ff0dff8",
        1893 => x"13860500",
        1894 => x"93050500",
        1895 => x"03a50186",
        1896 => x"6f004000",
        1897 => x"130101ff",
        1898 => x"23248100",
        1899 => x"23229100",
        1900 => x"13040500",
        1901 => x"13850500",
        1902 => x"93050600",
        1903 => x"23261100",
        1904 => x"23a20186",
        1905 => x"efe00fcc",
        1906 => x"9307f0ff",
        1907 => x"6318f500",
        1908 => x"83a74186",
        1909 => x"63840700",
        1910 => x"2320f400",
        1911 => x"8320c100",
        1912 => x"03248100",
        1913 => x"83244100",
        1914 => x"13010101",
        1915 => x"67800000",
        1916 => x"130101fe",
        1917 => x"23282101",
        1918 => x"03a98500",
        1919 => x"232c8100",
        1920 => x"23263101",
        1921 => x"23244101",
        1922 => x"23225101",
        1923 => x"232e1100",
        1924 => x"232a9100",
        1925 => x"23206101",
        1926 => x"83aa0500",
        1927 => x"13840500",
        1928 => x"130a0600",
        1929 => x"93890600",
        1930 => x"63ee2609",
        1931 => x"83d7c500",
        1932 => x"13f70748",
        1933 => x"63060708",
        1934 => x"83264401",
        1935 => x"83a50501",
        1936 => x"130b0500",
        1937 => x"13971600",
        1938 => x"3307d700",
        1939 => x"9354f701",
        1940 => x"b384e400",
        1941 => x"b38aba40",
        1942 => x"13871900",
        1943 => x"93d41440",
        1944 => x"33075701",
        1945 => x"63f4e400",
        1946 => x"93040700",
        1947 => x"93f70740",
        1948 => x"6386070a",
        1949 => x"93850400",
        1950 => x"13050b00",
        1951 => x"ef00d066",
        1952 => x"13090500",
        1953 => x"630c050a",
        1954 => x"83250401",
        1955 => x"13860a00",
        1956 => x"eff09fc5",
        1957 => x"8357c400",
        1958 => x"93f7f7b7",
        1959 => x"93e70708",
        1960 => x"2316f400",
        1961 => x"23282401",
        1962 => x"232a9400",
        1963 => x"33095901",
        1964 => x"b3845441",
        1965 => x"23202401",
        1966 => x"23249400",
        1967 => x"13890900",
        1968 => x"63f42901",
        1969 => x"13890900",
        1970 => x"03250400",
        1971 => x"13060900",
        1972 => x"93050a00",
        1973 => x"eff09fc3",
        1974 => x"83278400",
        1975 => x"13050000",
        1976 => x"b3872741",
        1977 => x"2324f400",
        1978 => x"83270400",
        1979 => x"b3872701",
        1980 => x"2320f400",
        1981 => x"8320c101",
        1982 => x"03248101",
        1983 => x"83244101",
        1984 => x"03290101",
        1985 => x"8329c100",
        1986 => x"032a8100",
        1987 => x"832a4100",
        1988 => x"032b0100",
        1989 => x"13010102",
        1990 => x"67800000",
        1991 => x"13860400",
        1992 => x"13050b00",
        1993 => x"ef005071",
        1994 => x"13090500",
        1995 => x"e31c05f6",
        1996 => x"83250401",
        1997 => x"13050b00",
        1998 => x"ef00904b",
        1999 => x"9307c000",
        2000 => x"2320fb00",
        2001 => x"8357c400",
        2002 => x"1305f0ff",
        2003 => x"93e70704",
        2004 => x"2316f400",
        2005 => x"6ff01ffa",
        2006 => x"83278600",
        2007 => x"130101fd",
        2008 => x"232e3101",
        2009 => x"23286101",
        2010 => x"23261102",
        2011 => x"23248102",
        2012 => x"23229102",
        2013 => x"23202103",
        2014 => x"232c4101",
        2015 => x"232a5101",
        2016 => x"23267101",
        2017 => x"23248101",
        2018 => x"032b0600",
        2019 => x"93090600",
        2020 => x"63980712",
        2021 => x"13050000",
        2022 => x"8320c102",
        2023 => x"03248102",
        2024 => x"23a20900",
        2025 => x"83244102",
        2026 => x"03290102",
        2027 => x"8329c101",
        2028 => x"032a8101",
        2029 => x"832a4101",
        2030 => x"032b0101",
        2031 => x"832bc100",
        2032 => x"032c8100",
        2033 => x"13010103",
        2034 => x"67800000",
        2035 => x"832a0b00",
        2036 => x"032c4b00",
        2037 => x"130b8b00",
        2038 => x"03298400",
        2039 => x"832b0400",
        2040 => x"e3060cfe",
        2041 => x"636a2c09",
        2042 => x"8357c400",
        2043 => x"13f70748",
        2044 => x"63040708",
        2045 => x"83264401",
        2046 => x"83250401",
        2047 => x"13971600",
        2048 => x"3307d700",
        2049 => x"9354f701",
        2050 => x"b38bbb40",
        2051 => x"b384e400",
        2052 => x"13871b00",
        2053 => x"93d41440",
        2054 => x"33078701",
        2055 => x"63f4e400",
        2056 => x"93040700",
        2057 => x"93f70740",
        2058 => x"6386070a",
        2059 => x"93850400",
        2060 => x"13050a00",
        2061 => x"ef00504b",
        2062 => x"13090500",
        2063 => x"630c050a",
        2064 => x"83250401",
        2065 => x"13860b00",
        2066 => x"eff01faa",
        2067 => x"8357c400",
        2068 => x"93f7f7b7",
        2069 => x"93e70708",
        2070 => x"2316f400",
        2071 => x"23282401",
        2072 => x"232a9400",
        2073 => x"33097901",
        2074 => x"b3847441",
        2075 => x"23202401",
        2076 => x"23249400",
        2077 => x"13090c00",
        2078 => x"63742c01",
        2079 => x"13090c00",
        2080 => x"03250400",
        2081 => x"93850a00",
        2082 => x"13060900",
        2083 => x"eff01fa8",
        2084 => x"83278400",
        2085 => x"b38a8a01",
        2086 => x"b3872741",
        2087 => x"2324f400",
        2088 => x"83270400",
        2089 => x"b3872701",
        2090 => x"2320f400",
        2091 => x"83a78900",
        2092 => x"b3878741",
        2093 => x"23a4f900",
        2094 => x"639a0700",
        2095 => x"6ff09fed",
        2096 => x"130a0500",
        2097 => x"13840500",
        2098 => x"930a0000",
        2099 => x"130c0000",
        2100 => x"6ff09ff0",
        2101 => x"13860400",
        2102 => x"13050a00",
        2103 => x"ef00d055",
        2104 => x"13090500",
        2105 => x"e31c05f6",
        2106 => x"83250401",
        2107 => x"13050a00",
        2108 => x"ef001030",
        2109 => x"9307c000",
        2110 => x"2320fa00",
        2111 => x"8357c400",
        2112 => x"1305f0ff",
        2113 => x"93e70704",
        2114 => x"2316f400",
        2115 => x"23a40900",
        2116 => x"6ff09fe8",
        2117 => x"83d7c500",
        2118 => x"130101f5",
        2119 => x"2324810a",
        2120 => x"2322910a",
        2121 => x"2320210b",
        2122 => x"232c4109",
        2123 => x"2326110a",
        2124 => x"232e3109",
        2125 => x"232a5109",
        2126 => x"23286109",
        2127 => x"23267109",
        2128 => x"23248109",
        2129 => x"23229109",
        2130 => x"2320a109",
        2131 => x"232eb107",
        2132 => x"93f70708",
        2133 => x"130a0500",
        2134 => x"13890500",
        2135 => x"93040600",
        2136 => x"13840600",
        2137 => x"63880706",
        2138 => x"83a70501",
        2139 => x"63940706",
        2140 => x"93050004",
        2141 => x"ef005037",
        2142 => x"2320a900",
        2143 => x"2328a900",
        2144 => x"63160504",
        2145 => x"9307c000",
        2146 => x"2320fa00",
        2147 => x"1305f0ff",
        2148 => x"8320c10a",
        2149 => x"0324810a",
        2150 => x"8324410a",
        2151 => x"0329010a",
        2152 => x"8329c109",
        2153 => x"032a8109",
        2154 => x"832a4109",
        2155 => x"032b0109",
        2156 => x"832bc108",
        2157 => x"032c8108",
        2158 => x"832c4108",
        2159 => x"032d0108",
        2160 => x"832dc107",
        2161 => x"1301010b",
        2162 => x"67800000",
        2163 => x"93070004",
        2164 => x"232af900",
        2165 => x"93070002",
        2166 => x"a304f102",
        2167 => x"93070003",
        2168 => x"23220102",
        2169 => x"2305f102",
        2170 => x"23268100",
        2171 => x"930c5002",
        2172 => x"373b0000",
        2173 => x"b73b0000",
        2174 => x"373d0000",
        2175 => x"372c0000",
        2176 => x"930a0000",
        2177 => x"13840400",
        2178 => x"83470400",
        2179 => x"63840700",
        2180 => x"6398970d",
        2181 => x"b30d9440",
        2182 => x"63069402",
        2183 => x"93860d00",
        2184 => x"13860400",
        2185 => x"93050900",
        2186 => x"13050a00",
        2187 => x"eff05fbc",
        2188 => x"9307f0ff",
        2189 => x"630af524",
        2190 => x"83274102",
        2191 => x"b387b701",
        2192 => x"2322f102",
        2193 => x"83470400",
        2194 => x"63800724",
        2195 => x"9307f0ff",
        2196 => x"93041400",
        2197 => x"23280100",
        2198 => x"232e0100",
        2199 => x"232af100",
        2200 => x"232c0100",
        2201 => x"a3090104",
        2202 => x"23240106",
        2203 => x"930d1000",
        2204 => x"83c50400",
        2205 => x"13065000",
        2206 => x"13054b28",
        2207 => x"ef001015",
        2208 => x"83270101",
        2209 => x"13841400",
        2210 => x"63100506",
        2211 => x"13f70701",
        2212 => x"63060700",
        2213 => x"13070002",
        2214 => x"a309e104",
        2215 => x"13f78700",
        2216 => x"63060700",
        2217 => x"1307b002",
        2218 => x"a309e104",
        2219 => x"83c60400",
        2220 => x"1307a002",
        2221 => x"6388e604",
        2222 => x"0327c101",
        2223 => x"13840400",
        2224 => x"93070000",
        2225 => x"13069000",
        2226 => x"83460400",
        2227 => x"93051400",
        2228 => x"938606fd",
        2229 => x"6376d610",
        2230 => x"63900704",
        2231 => x"6f004005",
        2232 => x"13041400",
        2233 => x"6ff05ff2",
        2234 => x"13074b28",
        2235 => x"3305e540",
        2236 => x"3395ad00",
        2237 => x"b3e7a700",
        2238 => x"2328f100",
        2239 => x"93040400",
        2240 => x"6ff01ff7",
        2241 => x"0327c100",
        2242 => x"93064700",
        2243 => x"03270700",
        2244 => x"2326d100",
        2245 => x"63460700",
        2246 => x"232ee100",
        2247 => x"6f004001",
        2248 => x"3307e040",
        2249 => x"93e72700",
        2250 => x"232ee100",
        2251 => x"2328f100",
        2252 => x"03470400",
        2253 => x"9307e002",
        2254 => x"6316f702",
        2255 => x"03471400",
        2256 => x"9307a002",
        2257 => x"6310f70c",
        2258 => x"8327c100",
        2259 => x"13042400",
        2260 => x"13874700",
        2261 => x"83a70700",
        2262 => x"2326e100",
        2263 => x"63c0070a",
        2264 => x"232af100",
        2265 => x"83450400",
        2266 => x"13063000",
        2267 => x"1385cb28",
        2268 => x"ef00d005",
        2269 => x"63020502",
        2270 => x"9387cb28",
        2271 => x"3305f540",
        2272 => x"83270101",
        2273 => x"13070004",
        2274 => x"3317a700",
        2275 => x"b3e7e700",
        2276 => x"13041400",
        2277 => x"2328f100",
        2278 => x"83450400",
        2279 => x"13066000",
        2280 => x"13050d29",
        2281 => x"93041400",
        2282 => x"2304b102",
        2283 => x"ef001002",
        2284 => x"6308050e",
        2285 => x"63960a0a",
        2286 => x"03270101",
        2287 => x"8327c100",
        2288 => x"13770710",
        2289 => x"63060708",
        2290 => x"93874700",
        2291 => x"2326f100",
        2292 => x"83274102",
        2293 => x"b3873701",
        2294 => x"2322f102",
        2295 => x"6ff09fe2",
        2296 => x"93172700",
        2297 => x"b387e700",
        2298 => x"93971700",
        2299 => x"3387d700",
        2300 => x"13840500",
        2301 => x"93071000",
        2302 => x"6ff01fed",
        2303 => x"9307f0ff",
        2304 => x"6ff01ff6",
        2305 => x"13041400",
        2306 => x"232a0100",
        2307 => x"93070000",
        2308 => x"13070000",
        2309 => x"13069000",
        2310 => x"83460400",
        2311 => x"93051400",
        2312 => x"938606fd",
        2313 => x"6378d600",
        2314 => x"e38e07f2",
        2315 => x"232ae100",
        2316 => x"6ff05ff3",
        2317 => x"93172700",
        2318 => x"b387e700",
        2319 => x"93971700",
        2320 => x"3387d700",
        2321 => x"13840500",
        2322 => x"93071000",
        2323 => x"6ff0dffc",
        2324 => x"93877700",
        2325 => x"93f787ff",
        2326 => x"93878700",
        2327 => x"6ff01ff7",
        2328 => x"1307c100",
        2329 => x"93060cdf",
        2330 => x"13060900",
        2331 => x"93050101",
        2332 => x"13050a00",
        2333 => x"97000000",
        2334 => x"e7000000",
        2335 => x"9307f0ff",
        2336 => x"93090500",
        2337 => x"e316f5f4",
        2338 => x"8357c900",
        2339 => x"1305f0ff",
        2340 => x"93f70704",
        2341 => x"e39e07ce",
        2342 => x"03254102",
        2343 => x"6ff05fcf",
        2344 => x"1307c100",
        2345 => x"93060cdf",
        2346 => x"13060900",
        2347 => x"93050101",
        2348 => x"13050a00",
        2349 => x"ef00801b",
        2350 => x"6ff05ffc",
        2351 => x"130101fd",
        2352 => x"232c4101",
        2353 => x"83a70501",
        2354 => x"130a0700",
        2355 => x"03a78500",
        2356 => x"23248102",
        2357 => x"23202103",
        2358 => x"232e3101",
        2359 => x"232a5101",
        2360 => x"23261102",
        2361 => x"23229102",
        2362 => x"23286101",
        2363 => x"23267101",
        2364 => x"93090500",
        2365 => x"13840500",
        2366 => x"13090600",
        2367 => x"938a0600",
        2368 => x"63d4e700",
        2369 => x"93070700",
        2370 => x"2320f900",
        2371 => x"03473404",
        2372 => x"63060700",
        2373 => x"93871700",
        2374 => x"2320f900",
        2375 => x"83270400",
        2376 => x"93f70702",
        2377 => x"63880700",
        2378 => x"83270900",
        2379 => x"93872700",
        2380 => x"2320f900",
        2381 => x"83240400",
        2382 => x"93f46400",
        2383 => x"639e0400",
        2384 => x"130b9401",
        2385 => x"930bf0ff",
        2386 => x"8327c400",
        2387 => x"03270900",
        2388 => x"b387e740",
        2389 => x"63c2f408",
        2390 => x"83473404",
        2391 => x"b336f000",
        2392 => x"83270400",
        2393 => x"93f70702",
        2394 => x"6390070c",
        2395 => x"13063404",
        2396 => x"93850a00",
        2397 => x"13850900",
        2398 => x"e7000a00",
        2399 => x"9307f0ff",
        2400 => x"6308f506",
        2401 => x"83270400",
        2402 => x"13074000",
        2403 => x"93040000",
        2404 => x"93f76700",
        2405 => x"639ce700",
        2406 => x"8324c400",
        2407 => x"83270900",
        2408 => x"b384f440",
        2409 => x"63d40400",
        2410 => x"93040000",
        2411 => x"83278400",
        2412 => x"03270401",
        2413 => x"6356f700",
        2414 => x"b387e740",
        2415 => x"b384f400",
        2416 => x"13090000",
        2417 => x"1304a401",
        2418 => x"130bf0ff",
        2419 => x"63902409",
        2420 => x"13050000",
        2421 => x"6f000002",
        2422 => x"93061000",
        2423 => x"13060b00",
        2424 => x"93850a00",
        2425 => x"13850900",
        2426 => x"e7000a00",
        2427 => x"631a7503",
        2428 => x"1305f0ff",
        2429 => x"8320c102",
        2430 => x"03248102",
        2431 => x"83244102",
        2432 => x"03290102",
        2433 => x"8329c101",
        2434 => x"032a8101",
        2435 => x"832a4101",
        2436 => x"032b0101",
        2437 => x"832bc100",
        2438 => x"13010103",
        2439 => x"67800000",
        2440 => x"93841400",
        2441 => x"6ff05ff2",
        2442 => x"3307d400",
        2443 => x"13060003",
        2444 => x"a301c704",
        2445 => x"03475404",
        2446 => x"93871600",
        2447 => x"b307f400",
        2448 => x"93862600",
        2449 => x"a381e704",
        2450 => x"6ff05ff2",
        2451 => x"93061000",
        2452 => x"13060400",
        2453 => x"93850a00",
        2454 => x"13850900",
        2455 => x"e7000a00",
        2456 => x"e30865f9",
        2457 => x"13091900",
        2458 => x"6ff05ff6",
        2459 => x"130101fc",
        2460 => x"232c8102",
        2461 => x"23244103",
        2462 => x"23225103",
        2463 => x"23206103",
        2464 => x"232e1102",
        2465 => x"232a9102",
        2466 => x"23282103",
        2467 => x"23263103",
        2468 => x"232e7101",
        2469 => x"232c8101",
        2470 => x"232a9101",
        2471 => x"83c78501",
        2472 => x"138b0600",
        2473 => x"93068007",
        2474 => x"130a0500",
        2475 => x"13840500",
        2476 => x"930a0600",
        2477 => x"63eef600",
        2478 => x"93062006",
        2479 => x"938b3504",
        2480 => x"63ecf600",
        2481 => x"6380072a",
        2482 => x"93068005",
        2483 => x"6388d724",
        2484 => x"930c2404",
        2485 => x"6f000004",
        2486 => x"1388d7f9",
        2487 => x"1378f80f",
        2488 => x"93065001",
        2489 => x"e3e606ff",
        2490 => x"b7360000",
        2491 => x"9386062c",
        2492 => x"13182800",
        2493 => x"3308d800",
        2494 => x"83260800",
        2495 => x"67800600",
        2496 => x"83270700",
        2497 => x"938c2504",
        2498 => x"93864700",
        2499 => x"83a70700",
        2500 => x"2320d700",
        2501 => x"2301f404",
        2502 => x"93071000",
        2503 => x"6f004028",
        2504 => x"83a70500",
        2505 => x"03260700",
        2506 => x"93f50708",
        2507 => x"93064600",
        2508 => x"63860502",
        2509 => x"83240600",
        2510 => x"2320d700",
        2511 => x"37390000",
        2512 => x"63d80400",
        2513 => x"9307d002",
        2514 => x"b3049040",
        2515 => x"a301f404",
        2516 => x"13098929",
        2517 => x"9309a000",
        2518 => x"6f00c00d",
        2519 => x"83240600",
        2520 => x"93f70704",
        2521 => x"2320d700",
        2522 => x"e38a07fc",
        2523 => x"93940401",
        2524 => x"93d40441",
        2525 => x"6ff09ffc",
        2526 => x"03a60500",
        2527 => x"83260700",
        2528 => x"13750608",
        2529 => x"93854600",
        2530 => x"63080500",
        2531 => x"2320b700",
        2532 => x"83a40600",
        2533 => x"6f004001",
        2534 => x"13760604",
        2535 => x"2320b700",
        2536 => x"e30806fe",
        2537 => x"83d40600",
        2538 => x"37390000",
        2539 => x"1307f006",
        2540 => x"13098929",
        2541 => x"9309a000",
        2542 => x"639ce706",
        2543 => x"93098000",
        2544 => x"6f000007",
        2545 => x"83a70500",
        2546 => x"93e70702",
        2547 => x"23a0f500",
        2548 => x"37390000",
        2549 => x"93078007",
        2550 => x"1309c92a",
        2551 => x"a302f404",
        2552 => x"83270400",
        2553 => x"83260700",
        2554 => x"13f60708",
        2555 => x"83a40600",
        2556 => x"93864600",
        2557 => x"631a0600",
        2558 => x"13f60704",
        2559 => x"63060600",
        2560 => x"93940401",
        2561 => x"93d40401",
        2562 => x"2320d700",
        2563 => x"13f71700",
        2564 => x"63060700",
        2565 => x"93e70702",
        2566 => x"2320f400",
        2567 => x"93090001",
        2568 => x"63980400",
        2569 => x"83270400",
        2570 => x"93f7f7fd",
        2571 => x"2320f400",
        2572 => x"a3010404",
        2573 => x"83274400",
        2574 => x"2324f400",
        2575 => x"63c80700",
        2576 => x"03270400",
        2577 => x"1377b7ff",
        2578 => x"2320e400",
        2579 => x"63960400",
        2580 => x"938c0b00",
        2581 => x"638e0702",
        2582 => x"938c0b00",
        2583 => x"93850900",
        2584 => x"13850400",
        2585 => x"eff04fa0",
        2586 => x"3305a900",
        2587 => x"83470500",
        2588 => x"93850900",
        2589 => x"13850400",
        2590 => x"a38ffcfe",
        2591 => x"138c0400",
        2592 => x"eff00f9a",
        2593 => x"938cfcff",
        2594 => x"93040500",
        2595 => x"e3783cfd",
        2596 => x"93078000",
        2597 => x"6394f902",
        2598 => x"83270400",
        2599 => x"93f71700",
        2600 => x"638e0700",
        2601 => x"03274400",
        2602 => x"83270401",
        2603 => x"63c8e700",
        2604 => x"93070003",
        2605 => x"a38ffcfe",
        2606 => x"938cfcff",
        2607 => x"b38b9b41",
        2608 => x"23287401",
        2609 => x"13070b00",
        2610 => x"93860a00",
        2611 => x"1306c100",
        2612 => x"93050400",
        2613 => x"13050a00",
        2614 => x"eff05fbe",
        2615 => x"9304f0ff",
        2616 => x"6316950c",
        2617 => x"1305f0ff",
        2618 => x"8320c103",
        2619 => x"03248103",
        2620 => x"83244103",
        2621 => x"03290103",
        2622 => x"8329c102",
        2623 => x"032a8102",
        2624 => x"832a4102",
        2625 => x"032b0102",
        2626 => x"832bc101",
        2627 => x"032c8101",
        2628 => x"832c4101",
        2629 => x"13010104",
        2630 => x"67800000",
        2631 => x"37390000",
        2632 => x"13098929",
        2633 => x"6ff09feb",
        2634 => x"83a60500",
        2635 => x"83270700",
        2636 => x"03a64501",
        2637 => x"13f50608",
        2638 => x"93854700",
        2639 => x"630a0500",
        2640 => x"2320b700",
        2641 => x"83a70700",
        2642 => x"23a0c700",
        2643 => x"6f008001",
        2644 => x"2320b700",
        2645 => x"93f60604",
        2646 => x"83a70700",
        2647 => x"e38606fe",
        2648 => x"2390c700",
        2649 => x"23280400",
        2650 => x"938c0b00",
        2651 => x"6ff09ff5",
        2652 => x"83270700",
        2653 => x"03a64500",
        2654 => x"93050000",
        2655 => x"93864700",
        2656 => x"2320d700",
        2657 => x"83ac0700",
        2658 => x"13850c00",
        2659 => x"ef000024",
        2660 => x"63060500",
        2661 => x"33059541",
        2662 => x"2322a400",
        2663 => x"83274400",
        2664 => x"2328f400",
        2665 => x"a3010404",
        2666 => x"6ff0dff1",
        2667 => x"83260401",
        2668 => x"13860c00",
        2669 => x"93850a00",
        2670 => x"13050a00",
        2671 => x"e7000b00",
        2672 => x"e30295f2",
        2673 => x"83270400",
        2674 => x"93f72700",
        2675 => x"63940704",
        2676 => x"8327c100",
        2677 => x"0325c400",
        2678 => x"e358f5f0",
        2679 => x"13850700",
        2680 => x"6ff09ff0",
        2681 => x"93061000",
        2682 => x"13060900",
        2683 => x"93850a00",
        2684 => x"13050a00",
        2685 => x"e7000b00",
        2686 => x"e30635ef",
        2687 => x"93841400",
        2688 => x"8327c400",
        2689 => x"0327c100",
        2690 => x"b387e740",
        2691 => x"e3ccf4fc",
        2692 => x"6ff01ffc",
        2693 => x"93040000",
        2694 => x"13099401",
        2695 => x"9309f0ff",
        2696 => x"6ff01ffe",
        2697 => x"130101ff",
        2698 => x"23248100",
        2699 => x"13840500",
        2700 => x"83a50500",
        2701 => x"23229100",
        2702 => x"23261100",
        2703 => x"93040500",
        2704 => x"63840500",
        2705 => x"eff01ffe",
        2706 => x"93050400",
        2707 => x"03248100",
        2708 => x"8320c100",
        2709 => x"13850400",
        2710 => x"83244100",
        2711 => x"13010101",
        2712 => x"6f000019",
        2713 => x"83a70186",
        2714 => x"6380a716",
        2715 => x"83274502",
        2716 => x"130101fe",
        2717 => x"232c8100",
        2718 => x"232e1100",
        2719 => x"232a9100",
        2720 => x"23282101",
        2721 => x"23263101",
        2722 => x"13040500",
        2723 => x"63840702",
        2724 => x"83a7c700",
        2725 => x"93040000",
        2726 => x"13090008",
        2727 => x"6392070e",
        2728 => x"83274402",
        2729 => x"83a50700",
        2730 => x"63860500",
        2731 => x"13050400",
        2732 => x"ef000014",
        2733 => x"83254401",
        2734 => x"63860500",
        2735 => x"13050400",
        2736 => x"ef000013",
        2737 => x"83254402",
        2738 => x"63860500",
        2739 => x"13050400",
        2740 => x"ef000012",
        2741 => x"83258403",
        2742 => x"63860500",
        2743 => x"13050400",
        2744 => x"ef000011",
        2745 => x"8325c403",
        2746 => x"63860500",
        2747 => x"13050400",
        2748 => x"ef000010",
        2749 => x"83250404",
        2750 => x"63860500",
        2751 => x"13050400",
        2752 => x"ef00000f",
        2753 => x"8325c405",
        2754 => x"63860500",
        2755 => x"13050400",
        2756 => x"ef00000e",
        2757 => x"83258405",
        2758 => x"63860500",
        2759 => x"13050400",
        2760 => x"ef00000d",
        2761 => x"83254403",
        2762 => x"63860500",
        2763 => x"13050400",
        2764 => x"ef00000c",
        2765 => x"83278401",
        2766 => x"638a0706",
        2767 => x"83278402",
        2768 => x"13050400",
        2769 => x"e7800700",
        2770 => x"83258404",
        2771 => x"63800506",
        2772 => x"13050400",
        2773 => x"03248101",
        2774 => x"8320c101",
        2775 => x"83244101",
        2776 => x"03290101",
        2777 => x"8329c100",
        2778 => x"13010102",
        2779 => x"6ff09feb",
        2780 => x"b3859500",
        2781 => x"83a50500",
        2782 => x"63900502",
        2783 => x"93844400",
        2784 => x"83274402",
        2785 => x"83a5c700",
        2786 => x"e39424ff",
        2787 => x"13050400",
        2788 => x"ef000006",
        2789 => x"6ff0dff0",
        2790 => x"83a90500",
        2791 => x"13050400",
        2792 => x"ef000005",
        2793 => x"93850900",
        2794 => x"6ff01ffd",
        2795 => x"8320c101",
        2796 => x"03248101",
        2797 => x"83244101",
        2798 => x"03290101",
        2799 => x"8329c100",
        2800 => x"13010102",
        2801 => x"67800000",
        2802 => x"67800000",
        2803 => x"93f5f50f",
        2804 => x"3306c500",
        2805 => x"6316c500",
        2806 => x"13050000",
        2807 => x"67800000",
        2808 => x"83470500",
        2809 => x"e38cb7fe",
        2810 => x"13051500",
        2811 => x"6ff09ffe",
        2812 => x"638a050e",
        2813 => x"83a7c5ff",
        2814 => x"130101fe",
        2815 => x"232c8100",
        2816 => x"232e1100",
        2817 => x"1384c5ff",
        2818 => x"63d40700",
        2819 => x"3304f400",
        2820 => x"2326a100",
        2821 => x"ef000034",
        2822 => x"83a78186",
        2823 => x"0325c100",
        2824 => x"639e0700",
        2825 => x"23220400",
        2826 => x"23a48186",
        2827 => x"03248101",
        2828 => x"8320c101",
        2829 => x"13010102",
        2830 => x"6f000032",
        2831 => x"6374f402",
        2832 => x"03260400",
        2833 => x"b306c400",
        2834 => x"639ad700",
        2835 => x"83a60700",
        2836 => x"83a74700",
        2837 => x"b386c600",
        2838 => x"2320d400",
        2839 => x"2322f400",
        2840 => x"6ff09ffc",
        2841 => x"13870700",
        2842 => x"83a74700",
        2843 => x"63840700",
        2844 => x"e37af4fe",
        2845 => x"83260700",
        2846 => x"3306d700",
        2847 => x"63188602",
        2848 => x"03260400",
        2849 => x"b386c600",
        2850 => x"2320d700",
        2851 => x"3306d700",
        2852 => x"e39ec7f8",
        2853 => x"03a60700",
        2854 => x"83a74700",
        2855 => x"b306d600",
        2856 => x"2320d700",
        2857 => x"2322f700",
        2858 => x"6ff05ff8",
        2859 => x"6378c400",
        2860 => x"9307c000",
        2861 => x"2320f500",
        2862 => x"6ff05ff7",
        2863 => x"03260400",
        2864 => x"b306c400",
        2865 => x"639ad700",
        2866 => x"83a60700",
        2867 => x"83a74700",
        2868 => x"b386c600",
        2869 => x"2320d400",
        2870 => x"2322f400",
        2871 => x"23228700",
        2872 => x"6ff0dff4",
        2873 => x"67800000",
        2874 => x"130101fe",
        2875 => x"232a9100",
        2876 => x"93843500",
        2877 => x"93f4c4ff",
        2878 => x"23282101",
        2879 => x"232e1100",
        2880 => x"232c8100",
        2881 => x"23263101",
        2882 => x"93848400",
        2883 => x"9307c000",
        2884 => x"13090500",
        2885 => x"63f4f406",
        2886 => x"9304c000",
        2887 => x"63e2b406",
        2888 => x"13050900",
        2889 => x"ef000023",
        2890 => x"03a78186",
        2891 => x"93868186",
        2892 => x"13040700",
        2893 => x"631a0406",
        2894 => x"1384c186",
        2895 => x"83270400",
        2896 => x"639a0700",
        2897 => x"93050000",
        2898 => x"13050900",
        2899 => x"ef00001c",
        2900 => x"2320a400",
        2901 => x"93850400",
        2902 => x"13050900",
        2903 => x"ef00001b",
        2904 => x"9309f0ff",
        2905 => x"631a350b",
        2906 => x"9307c000",
        2907 => x"2320f900",
        2908 => x"13050900",
        2909 => x"ef00401e",
        2910 => x"6f000001",
        2911 => x"e3d004fa",
        2912 => x"9307c000",
        2913 => x"2320f900",
        2914 => x"13050000",
        2915 => x"8320c101",
        2916 => x"03248101",
        2917 => x"83244101",
        2918 => x"03290101",
        2919 => x"8329c100",
        2920 => x"13010102",
        2921 => x"67800000",
        2922 => x"83270400",
        2923 => x"b3879740",
        2924 => x"63ce0704",
        2925 => x"1306b000",
        2926 => x"637af600",
        2927 => x"2320f400",
        2928 => x"3304f400",
        2929 => x"23209400",
        2930 => x"6f000001",
        2931 => x"83274400",
        2932 => x"631a8702",
        2933 => x"23a0f600",
        2934 => x"13050900",
        2935 => x"ef00c017",
        2936 => x"1305b400",
        2937 => x"93074400",
        2938 => x"137585ff",
        2939 => x"3307f540",
        2940 => x"e30ef5f8",
        2941 => x"3304e400",
        2942 => x"b387a740",
        2943 => x"2320f400",
        2944 => x"6ff0dff8",
        2945 => x"2322f700",
        2946 => x"6ff01ffd",
        2947 => x"13070400",
        2948 => x"03244400",
        2949 => x"6ff01ff2",
        2950 => x"13043500",
        2951 => x"1374c4ff",
        2952 => x"e30285fa",
        2953 => x"b305a440",
        2954 => x"13050900",
        2955 => x"ef00000e",
        2956 => x"e31a35f9",
        2957 => x"6ff05ff3",
        2958 => x"130101fe",
        2959 => x"232c8100",
        2960 => x"232e1100",
        2961 => x"232a9100",
        2962 => x"23282101",
        2963 => x"23263101",
        2964 => x"23244101",
        2965 => x"13040600",
        2966 => x"63940502",
        2967 => x"03248101",
        2968 => x"8320c101",
        2969 => x"83244101",
        2970 => x"03290101",
        2971 => x"8329c100",
        2972 => x"032a8100",
        2973 => x"93050600",
        2974 => x"13010102",
        2975 => x"6ff0dfe6",
        2976 => x"63180602",
        2977 => x"eff0dfd6",
        2978 => x"93040000",
        2979 => x"8320c101",
        2980 => x"03248101",
        2981 => x"03290101",
        2982 => x"8329c100",
        2983 => x"032a8100",
        2984 => x"13850400",
        2985 => x"83244101",
        2986 => x"13010102",
        2987 => x"67800000",
        2988 => x"130a0500",
        2989 => x"13890500",
        2990 => x"ef00400a",
        2991 => x"93090500",
        2992 => x"63688500",
        2993 => x"93571500",
        2994 => x"93040900",
        2995 => x"e3e087fc",
        2996 => x"93050400",
        2997 => x"13050a00",
        2998 => x"eff01fe1",
        2999 => x"93040500",
        3000 => x"e30605fa",
        3001 => x"13060400",
        3002 => x"63f48900",
        3003 => x"13860900",
        3004 => x"93050900",
        3005 => x"13850400",
        3006 => x"efe01fbf",
        3007 => x"93050900",
        3008 => x"13050a00",
        3009 => x"eff0dfce",
        3010 => x"6ff05ff8",
        3011 => x"130101ff",
        3012 => x"23248100",
        3013 => x"23229100",
        3014 => x"13040500",
        3015 => x"13850500",
        3016 => x"23261100",
        3017 => x"23a20186",
        3018 => x"efd08fc7",
        3019 => x"9307f0ff",
        3020 => x"6318f500",
        3021 => x"83a74186",
        3022 => x"63840700",
        3023 => x"2320f400",
        3024 => x"8320c100",
        3025 => x"03248100",
        3026 => x"83244100",
        3027 => x"13010101",
        3028 => x"67800000",
        3029 => x"67800000",
        3030 => x"67800000",
        3031 => x"83a7c5ff",
        3032 => x"1385c7ff",
        3033 => x"63d80700",
        3034 => x"b385a500",
        3035 => x"83a70500",
        3036 => x"3305f500",
        3037 => x"67800000",
        3038 => x"9308d005",
        3039 => x"73000000",
        3040 => x"63520502",
        3041 => x"130101ff",
        3042 => x"23248100",
        3043 => x"13040500",
        3044 => x"23261100",
        3045 => x"33048040",
        3046 => x"efe01fbb",
        3047 => x"23208500",
        3048 => x"6f000000",
        3049 => x"6f000000",
        3050 => x"10000000",
        3051 => x"00000000",
        3052 => x"037a5200",
        3053 => x"017c0101",
        3054 => x"1b0d0200",
        3055 => x"4c000000",
        3056 => x"18000000",
        3057 => x"78d4ffff",
        3058 => x"10060000",
        3059 => x"00440e30",
        3060 => x"70890394",
        3061 => x"06810188",
        3062 => x"02920493",
        3063 => x"05950796",
        3064 => x"08970998",
        3065 => x"0a990b9a",
        3066 => x"0c03a402",
        3067 => x"0ac144c8",
        3068 => x"44c944d2",
        3069 => x"44d344d4",
        3070 => x"44d544d6",
        3071 => x"44d744d8",
        3072 => x"44d944da",
        3073 => x"440e0044",
        3074 => x"0b000000",
        3075 => x"10000000",
        3076 => x"00000000",
        3077 => x"037a5200",
        3078 => x"017c0101",
        3079 => x"1b0d0200",
        3080 => x"50000000",
        3081 => x"18000000",
        3082 => x"24daffff",
        3083 => x"18050000",
        3084 => x"00440e40",
        3085 => x"74890381",
        3086 => x"01880292",
        3087 => x"04930594",
        3088 => x"06950796",
        3089 => x"08970998",
        3090 => x"0a990b9a",
        3091 => x"0c9b0d03",
        3092 => x"50010ac1",
        3093 => x"44c844c9",
        3094 => x"44d244d3",
        3095 => x"44d444d5",
        3096 => x"44d644d7",
        3097 => x"44d844d9",
        3098 => x"44da44db",
        3099 => x"440e0044",
        3100 => x"0b000000",
        3101 => x"10000000",
        3102 => x"00000000",
        3103 => x"037a5200",
        3104 => x"017c0101",
        3105 => x"1b0d0200",
        3106 => x"48000000",
        3107 => x"18000000",
        3108 => x"d4deffff",
        3109 => x"c0050000",
        3110 => x"00440e30",
        3111 => x"6c930581",
        3112 => x"01880289",
        3113 => x"03920494",
        3114 => x"06950796",
        3115 => x"08970998",
        3116 => x"0a990b03",
        3117 => x"54020ac1",
        3118 => x"44c844c9",
        3119 => x"44d344d4",
        3120 => x"44d544d6",
        3121 => x"44d744d8",
        3122 => x"44d94cd2",
        3123 => x"440e0044",
        3124 => x"0b000000",
        3125 => x"10000000",
        3126 => x"00000000",
        3127 => x"037a5200",
        3128 => x"017c0101",
        3129 => x"1b0d0200",
        3130 => x"4c000000",
        3131 => x"18000000",
        3132 => x"34e4ffff",
        3133 => x"d0040000",
        3134 => x"00440e30",
        3135 => x"70880289",
        3136 => x"03810192",
        3137 => x"04930594",
        3138 => x"06950796",
        3139 => x"08970998",
        3140 => x"0a990b9a",
        3141 => x"0c030c01",
        3142 => x"0ac144c8",
        3143 => x"44c944d2",
        3144 => x"44d344d4",
        3145 => x"44d544d6",
        3146 => x"44d744d8",
        3147 => x"44d944da",
        3148 => x"440e0044",
        3149 => x"0b000000",
        3150 => x"0d0a0d0a",
        3151 => x"54696d65",
        3152 => x"2073696e",
        3153 => x"6365206c",
        3154 => x"61737420",
        3155 => x"72657365",
        3156 => x"743a0d0a",
        3157 => x"00000000",
        3158 => x"256c642c",
        3159 => x"2530366c",
        3160 => x"64207c20",
        3161 => x"2530336c",
        3162 => x"643a2530",
        3163 => x"326c643a",
        3164 => x"2530326c",
        3165 => x"64202020",
        3166 => x"20202020",
        3167 => x"20202020",
        3168 => x"0d000000",
        3169 => x"00010202",
        3170 => x"03030303",
        3171 => x"04040404",
        3172 => x"04040404",
        3173 => x"05050505",
        3174 => x"05050505",
        3175 => x"05050505",
        3176 => x"05050505",
        3177 => x"06060606",
        3178 => x"06060606",
        3179 => x"06060606",
        3180 => x"06060606",
        3181 => x"06060606",
        3182 => x"06060606",
        3183 => x"06060606",
        3184 => x"06060606",
        3185 => x"07070707",
        3186 => x"07070707",
        3187 => x"07070707",
        3188 => x"07070707",
        3189 => x"07070707",
        3190 => x"07070707",
        3191 => x"07070707",
        3192 => x"07070707",
        3193 => x"07070707",
        3194 => x"07070707",
        3195 => x"07070707",
        3196 => x"07070707",
        3197 => x"07070707",
        3198 => x"07070707",
        3199 => x"07070707",
        3200 => x"07070707",
        3201 => x"08080808",
        3202 => x"08080808",
        3203 => x"08080808",
        3204 => x"08080808",
        3205 => x"08080808",
        3206 => x"08080808",
        3207 => x"08080808",
        3208 => x"08080808",
        3209 => x"08080808",
        3210 => x"08080808",
        3211 => x"08080808",
        3212 => x"08080808",
        3213 => x"08080808",
        3214 => x"08080808",
        3215 => x"08080808",
        3216 => x"08080808",
        3217 => x"08080808",
        3218 => x"08080808",
        3219 => x"08080808",
        3220 => x"08080808",
        3221 => x"08080808",
        3222 => x"08080808",
        3223 => x"08080808",
        3224 => x"08080808",
        3225 => x"08080808",
        3226 => x"08080808",
        3227 => x"08080808",
        3228 => x"08080808",
        3229 => x"08080808",
        3230 => x"08080808",
        3231 => x"08080808",
        3232 => x"08080808",
        3233 => x"232d302b",
        3234 => x"20000000",
        3235 => x"686c4c00",
        3236 => x"65666745",
        3237 => x"46470000",
        3238 => x"30313233",
        3239 => x"34353637",
        3240 => x"38394142",
        3241 => x"43444546",
        3242 => x"00000000",
        3243 => x"30313233",
        3244 => x"34353637",
        3245 => x"38396162",
        3246 => x"63646566",
        3247 => x"00000000",
        3248 => x"00270000",
        3249 => x"20270000",
        3250 => x"d0260000",
        3251 => x"d0260000",
        3252 => x"d0260000",
        3253 => x"d0260000",
        3254 => x"20270000",
        3255 => x"d0260000",
        3256 => x"d0260000",
        3257 => x"d0260000",
        3258 => x"d0260000",
        3259 => x"28290000",
        3260 => x"78270000",
        3261 => x"c4270000",
        3262 => x"d0260000",
        3263 => x"d0260000",
        3264 => x"70290000",
        3265 => x"d0260000",
        3266 => x"78270000",
        3267 => x"d0260000",
        3268 => x"d0260000",
        3269 => x"d0270000",
        3270 => x"00000020",
        3271 => x"00000000",
        3272 => x"00000000",
        3273 => x"00000000",
        3274 => x"00000000",
        3275 => x"00000000",
        3276 => x"00000000",
        3277 => x"00000000",
        3278 => x"00000000",
        3279 => x"00000000",
        3280 => x"00000000",
        3281 => x"00000000",
        3282 => x"00000000",
        3283 => x"00000000",
        3284 => x"00000000",
        3285 => x"00000000",
        3286 => x"00000000",
        3287 => x"00000000",
        3288 => x"00000000",
        3289 => x"00000000",
        3290 => x"00000000",
        3291 => x"00000000",
        3292 => x"00000000",
        3293 => x"00000000",
        3294 => x"00000000",
        3295 => x"00000020",
        others => (others => '-')
    );
end package processor_common_rom;
