-- srec2vhdl table generator
-- for input file string.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97",    1 => x"11",    2 => x"00",    3 => x"20", 
           4 => x"93",    5 => x"81",    6 => x"01",    7 => x"87", 
           8 => x"17",    9 => x"41",   10 => x"00",   11 => x"20", 
          12 => x"13",   13 => x"01",   14 => x"81",   15 => x"ff", 
          16 => x"33",   17 => x"04",   18 => x"01",   19 => x"00", 
          20 => x"b7",   21 => x"07",   22 => x"00",   23 => x"20", 
          24 => x"93",   25 => x"80",   26 => x"47",   27 => x"06", 
          28 => x"b7",   29 => x"07",   30 => x"00",   31 => x"20", 
          32 => x"93",   33 => x"84",   34 => x"47",   35 => x"06", 
          36 => x"13",   37 => x"09",   38 => x"40",   39 => x"29", 
          40 => x"6f",   41 => x"00",   42 => x"40",   43 => x"01", 
          44 => x"23",   45 => x"a0",   46 => x"00",   47 => x"00", 
          48 => x"93",   49 => x"87",   50 => x"00",   51 => x"00", 
          52 => x"93",   53 => x"80",   54 => x"47",   55 => x"00", 
          56 => x"83",   57 => x"a7",   58 => x"07",   59 => x"00", 
          60 => x"e3",   61 => x"e8",   62 => x"90",   63 => x"fe", 
          64 => x"b7",   65 => x"07",   66 => x"00",   67 => x"20", 
          68 => x"93",   69 => x"80",   70 => x"07",   71 => x"00", 
          72 => x"b7",   73 => x"07",   74 => x"00",   75 => x"20", 
          76 => x"93",   77 => x"84",   78 => x"07",   79 => x"06", 
          80 => x"6f",   81 => x"00",   82 => x"40",   83 => x"01", 
          84 => x"83",   85 => x"27",   86 => x"09",   87 => x"00", 
          88 => x"23",   89 => x"a0",   90 => x"f0",   91 => x"00", 
          92 => x"93",   93 => x"80",   94 => x"40",   95 => x"00", 
          96 => x"13",   97 => x"09",   98 => x"49",   99 => x"00", 
         100 => x"e3",  101 => x"e8",  102 => x"90",  103 => x"fe", 
         104 => x"ef",  105 => x"00",  106 => x"80",  107 => x"10", 
         108 => x"ef",  109 => x"00",  110 => x"c0",  111 => x"00", 
         112 => x"13",  113 => x"05",  114 => x"00",  115 => x"00", 
         116 => x"ef",  117 => x"00",  118 => x"00",  119 => x"0c", 
         120 => x"13",  121 => x"01",  122 => x"01",  123 => x"f7", 
         124 => x"23",  125 => x"26",  126 => x"11",  127 => x"08", 
         128 => x"23",  129 => x"24",  130 => x"81",  131 => x"08", 
         132 => x"13",  133 => x"04",  134 => x"01",  135 => x"09", 
         136 => x"93",  137 => x"07",  138 => x"80",  139 => x"27", 
         140 => x"03",  141 => x"a5",  142 => x"07",  143 => x"00", 
         144 => x"83",  145 => x"a5",  146 => x"47",  147 => x"00", 
         148 => x"03",  149 => x"a6",  150 => x"87",  151 => x"00", 
         152 => x"83",  153 => x"a6",  154 => x"c7",  155 => x"00", 
         156 => x"03",  157 => x"a7",  158 => x"07",  159 => x"01", 
         160 => x"83",  161 => x"a7",  162 => x"47",  163 => x"01", 
         164 => x"23",  165 => x"2c",  166 => x"a4",  167 => x"fc", 
         168 => x"23",  169 => x"2e",  170 => x"b4",  171 => x"fc", 
         172 => x"23",  173 => x"20",  174 => x"c4",  175 => x"fe", 
         176 => x"23",  177 => x"22",  178 => x"d4",  179 => x"fe", 
         180 => x"23",  181 => x"24",  182 => x"e4",  183 => x"fe", 
         184 => x"23",  185 => x"26",  186 => x"f4",  187 => x"fe", 
         188 => x"93",  189 => x"07",  190 => x"84",  191 => x"fd", 
         192 => x"13",  193 => x"85",  194 => x"07",  195 => x"00", 
         196 => x"ef",  197 => x"00",  198 => x"40",  199 => x"15", 
         200 => x"93",  201 => x"07",  202 => x"05",  203 => x"00", 
         204 => x"23",  205 => x"28",  206 => x"f4",  207 => x"f6", 
         208 => x"13",  209 => x"07",  210 => x"84",  211 => x"fd", 
         212 => x"93",  213 => x"07",  214 => x"44",  215 => x"f7", 
         216 => x"93",  217 => x"05",  218 => x"07",  219 => x"00", 
         220 => x"13",  221 => x"85",  222 => x"07",  223 => x"00", 
         224 => x"ef",  225 => x"00",  226 => x"c0",  227 => x"11", 
         228 => x"93",  229 => x"07",  230 => x"84",  231 => x"fd", 
         232 => x"93",  233 => x"85",  234 => x"07",  235 => x"00", 
         236 => x"13",  237 => x"05",  238 => x"00",  239 => x"27", 
         240 => x"ef",  241 => x"00",  242 => x"40",  243 => x"02", 
         244 => x"93",  245 => x"07",  246 => x"05",  247 => x"00", 
         248 => x"23",  249 => x"28",  250 => x"f4",  251 => x"f6", 
         252 => x"83",  253 => x"27",  254 => x"04",  255 => x"f7", 
         256 => x"13",  257 => x"85",  258 => x"07",  259 => x"00", 
         260 => x"83",  261 => x"20",  262 => x"c1",  263 => x"08", 
         264 => x"03",  265 => x"24",  266 => x"81",  267 => x"08", 
         268 => x"13",  269 => x"01",  270 => x"01",  271 => x"09", 
         272 => x"67",  273 => x"80",  274 => x"00",  275 => x"00", 
         276 => x"03",  277 => x"46",  278 => x"05",  279 => x"00", 
         280 => x"83",  281 => x"c6",  282 => x"05",  283 => x"00", 
         284 => x"13",  285 => x"05",  286 => x"15",  287 => x"00", 
         288 => x"93",  289 => x"85",  290 => x"15",  291 => x"00", 
         292 => x"63",  293 => x"14",  294 => x"d6",  295 => x"00", 
         296 => x"e3",  297 => x"16",  298 => x"06",  299 => x"fe", 
         300 => x"33",  301 => x"05",  302 => x"d6",  303 => x"40", 
         304 => x"67",  305 => x"80",  306 => x"00",  307 => x"00", 
         308 => x"13",  309 => x"01",  310 => x"01",  311 => x"ff", 
         312 => x"23",  313 => x"24",  314 => x"81",  315 => x"00", 
         316 => x"23",  317 => x"26",  318 => x"11",  319 => x"00", 
         320 => x"93",  321 => x"07",  322 => x"00",  323 => x"00", 
         324 => x"13",  325 => x"04",  326 => x"05",  327 => x"00", 
         328 => x"63",  329 => x"88",  330 => x"07",  331 => x"00", 
         332 => x"93",  333 => x"05",  334 => x"00",  335 => x"00", 
         336 => x"97",  337 => x"00",  338 => x"00",  339 => x"00", 
         340 => x"e7",  341 => x"00",  342 => x"00",  343 => x"00", 
         344 => x"03",  345 => x"25",  346 => x"00",  347 => x"29", 
         348 => x"83",  349 => x"27",  350 => x"85",  351 => x"02", 
         352 => x"63",  353 => x"84",  354 => x"07",  355 => x"00", 
         356 => x"e7",  357 => x"80",  358 => x"07",  359 => x"00", 
         360 => x"13",  361 => x"05",  362 => x"04",  363 => x"00", 
         364 => x"ef",  365 => x"00",  366 => x"80",  367 => x"0c", 
         368 => x"13",  369 => x"01",  370 => x"01",  371 => x"ff", 
         372 => x"23",  373 => x"24",  374 => x"81",  375 => x"00", 
         376 => x"23",  377 => x"22",  378 => x"91",  379 => x"00", 
         380 => x"93",  381 => x"07",  382 => x"40",  383 => x"29", 
         384 => x"13",  385 => x"04",  386 => x"40",  387 => x"29", 
         388 => x"33",  389 => x"04",  390 => x"f4",  391 => x"40", 
         392 => x"23",  393 => x"20",  394 => x"21",  395 => x"01", 
         396 => x"23",  397 => x"26",  398 => x"11",  399 => x"00", 
         400 => x"13",  401 => x"54",  402 => x"24",  403 => x"40", 
         404 => x"93",  405 => x"04",  406 => x"40",  407 => x"29", 
         408 => x"13",  409 => x"09",  410 => x"00",  411 => x"00", 
         412 => x"63",  413 => x"1c",  414 => x"89",  415 => x"02", 
         416 => x"93",  417 => x"07",  418 => x"40",  419 => x"29", 
         420 => x"13",  421 => x"04",  422 => x"40",  423 => x"29", 
         424 => x"33",  425 => x"04",  426 => x"f4",  427 => x"40", 
         428 => x"13",  429 => x"54",  430 => x"24",  431 => x"40", 
         432 => x"93",  433 => x"04",  434 => x"40",  435 => x"29", 
         436 => x"13",  437 => x"09",  438 => x"00",  439 => x"00", 
         440 => x"63",  441 => x"18",  442 => x"89",  443 => x"02", 
         444 => x"83",  445 => x"20",  446 => x"c1",  447 => x"00", 
         448 => x"03",  449 => x"24",  450 => x"81",  451 => x"00", 
         452 => x"83",  453 => x"24",  454 => x"41",  455 => x"00", 
         456 => x"03",  457 => x"29",  458 => x"01",  459 => x"00", 
         460 => x"13",  461 => x"01",  462 => x"01",  463 => x"01", 
         464 => x"67",  465 => x"80",  466 => x"00",  467 => x"00", 
         468 => x"83",  469 => x"a7",  470 => x"04",  471 => x"00", 
         472 => x"13",  473 => x"09",  474 => x"19",  475 => x"00", 
         476 => x"93",  477 => x"84",  478 => x"44",  479 => x"00", 
         480 => x"e7",  481 => x"80",  482 => x"07",  483 => x"00", 
         484 => x"6f",  485 => x"f0",  486 => x"9f",  487 => x"fb", 
         488 => x"83",  489 => x"a7",  490 => x"04",  491 => x"00", 
         492 => x"13",  493 => x"09",  494 => x"19",  495 => x"00", 
         496 => x"93",  497 => x"84",  498 => x"44",  499 => x"00", 
         500 => x"e7",  501 => x"80",  502 => x"07",  503 => x"00", 
         504 => x"6f",  505 => x"f0",  506 => x"1f",  507 => x"fc", 
         508 => x"93",  509 => x"07",  510 => x"05",  511 => x"00", 
         512 => x"03",  513 => x"c7",  514 => x"05",  515 => x"00", 
         516 => x"93",  517 => x"87",  518 => x"17",  519 => x"00", 
         520 => x"93",  521 => x"85",  522 => x"15",  523 => x"00", 
         524 => x"a3",  525 => x"8f",  526 => x"e7",  527 => x"fe", 
         528 => x"e3",  529 => x"18",  530 => x"07",  531 => x"fe", 
         532 => x"67",  533 => x"80",  534 => x"00",  535 => x"00", 
         536 => x"93",  537 => x"07",  538 => x"05",  539 => x"00", 
         540 => x"03",  541 => x"c7",  542 => x"07",  543 => x"00", 
         544 => x"93",  545 => x"87",  546 => x"17",  547 => x"00", 
         548 => x"e3",  549 => x"1c",  550 => x"07",  551 => x"fe", 
         552 => x"33",  553 => x"85",  554 => x"a7",  555 => x"40", 
         556 => x"13",  557 => x"05",  558 => x"f5",  559 => x"ff", 
         560 => x"67",  561 => x"80",  562 => x"00",  563 => x"00", 
         564 => x"93",  565 => x"08",  566 => x"d0",  567 => x"05", 
         568 => x"73",  569 => x"00",  570 => x"00",  571 => x"00", 
         572 => x"63",  573 => x"52",  574 => x"05",  575 => x"02", 
         576 => x"13",  577 => x"01",  578 => x"01",  579 => x"ff", 
         580 => x"23",  581 => x"24",  582 => x"81",  583 => x"00", 
         584 => x"13",  585 => x"04",  586 => x"05",  587 => x"00", 
         588 => x"23",  589 => x"26",  590 => x"11",  591 => x"00", 
         592 => x"33",  593 => x"04",  594 => x"80",  595 => x"40", 
         596 => x"ef",  597 => x"00",  598 => x"00",  599 => x"01", 
         600 => x"23",  601 => x"20",  602 => x"85",  603 => x"00", 
         604 => x"6f",  605 => x"00",  606 => x"00",  607 => x"00", 
         608 => x"6f",  609 => x"00",  610 => x"00",  611 => x"00", 
         612 => x"b7",  613 => x"07",  614 => x"00",  615 => x"20", 
         616 => x"03",  617 => x"a5",  618 => x"07",  619 => x"06", 
         620 => x"67",  621 => x"80",  622 => x"00",  623 => x"00", 
         624 => x"48",  625 => x"65",  626 => x"6c",  627 => x"6c", 
         628 => x"6f",  629 => x"00",  630 => x"00",  631 => x"00", 
         632 => x"48",  633 => x"65",  634 => x"6c",  635 => x"6c", 
         636 => x"6f",  637 => x"20",  638 => x"64",  639 => x"69", 
         640 => x"74",  641 => x"20",  642 => x"69",  643 => x"73", 
         644 => x"20",  645 => x"65",  646 => x"65",  647 => x"6e", 
         648 => x"20",  649 => x"73",  650 => x"74",  651 => x"72", 
         652 => x"69",  653 => x"6e",  654 => x"67",  655 => x"00", 
         656 => x"00",  657 => x"00",  658 => x"00",  659 => x"20", 
         660 => x"00",  661 => x"00",  662 => x"00",  663 => x"00", 
         664 => x"00",  665 => x"00",  666 => x"00",  667 => x"00", 
         668 => x"00",  669 => x"00",  670 => x"00",  671 => x"00", 
         672 => x"00",  673 => x"00",  674 => x"00",  675 => x"00", 
         676 => x"00",  677 => x"00",  678 => x"00",  679 => x"00", 
         680 => x"00",  681 => x"00",  682 => x"00",  683 => x"00", 
         684 => x"00",  685 => x"00",  686 => x"00",  687 => x"00", 
         688 => x"00",  689 => x"00",  690 => x"00",  691 => x"00", 
         692 => x"00",  693 => x"00",  694 => x"00",  695 => x"00", 
         696 => x"00",  697 => x"00",  698 => x"00",  699 => x"00", 
         700 => x"00",  701 => x"00",  702 => x"00",  703 => x"00", 
         704 => x"00",  705 => x"00",  706 => x"00",  707 => x"00", 
         708 => x"00",  709 => x"00",  710 => x"00",  711 => x"00", 
         712 => x"00",  713 => x"00",  714 => x"00",  715 => x"00", 
         716 => x"00",  717 => x"00",  718 => x"00",  719 => x"00", 
         720 => x"00",  721 => x"00",  722 => x"00",  723 => x"00", 
         724 => x"00",  725 => x"00",  726 => x"00",  727 => x"00", 
         728 => x"00",  729 => x"00",  730 => x"00",  731 => x"00", 
         732 => x"00",  733 => x"00",  734 => x"00",  735 => x"00", 
         736 => x"00",  737 => x"00",  738 => x"00",  739 => x"00", 
         740 => x"00",  741 => x"00",  742 => x"00",  743 => x"00", 
         744 => x"00",  745 => x"00",  746 => x"00",  747 => x"00", 
         748 => x"00",  749 => x"00",  750 => x"00",  751 => x"00", 
         752 => x"00",  753 => x"00",  754 => x"00",  755 => x"00", 
         756 => x"00",  757 => x"00",  758 => x"00",  759 => x"20", 
        others => (others => '-')
    );
end package processor_common_rom;
